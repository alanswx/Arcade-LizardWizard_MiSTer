library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"F1",X"4F",X"C3",X"59",X"00",X"21",X"16",X"40",X"11",X"17",X"40",X"01",X"08",X"00",X"36",
		X"40",X"ED",X"B0",X"3A",X"A1",X"4D",X"FE",X"00",X"C8",X"47",X"3E",X"3A",X"21",X"1D",X"40",X"77",
		X"2B",X"10",X"FC",X"C9",X"00",X"08",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"08",X"0A",X"21",X"02",X"40",X"11",X"03",
		X"40",X"01",X"08",X"00",X"36",X"40",X"ED",X"B0",X"3A",X"A2",X"4D",X"FE",X"00",X"C8",X"47",X"3E",
		X"3A",X"21",X"02",X"40",X"77",X"23",X"10",X"FC",X"C9",X"AF",X"06",X"08",X"21",X"00",X"50",X"77",
		X"23",X"10",X"FC",X"3A",X"00",X"50",X"CB",X"67",X"C2",X"57",X"03",X"AF",X"06",X"08",X"21",X"00",
		X"50",X"77",X"23",X"10",X"FC",X"C3",X"95",X"00",X"06",X"03",X"0E",X"0F",X"3E",X"21",X"ED",X"A0",
		X"CD",X"52",X"16",X"10",X"F7",X"23",X"23",X"3E",X"40",X"CD",X"52",X"16",X"CD",X"9C",X"11",X"3E",
		X"04",X"CD",X"E3",X"15",X"C9",X"3E",X"00",X"32",X"03",X"50",X"31",X"F1",X"4F",X"CD",X"24",X"12",
		X"F3",X"08",X"AF",X"08",X"21",X"00",X"40",X"CD",X"D2",X"02",X"08",X"CB",X"47",X"28",X"02",X"CB",
		X"D7",X"CB",X"4F",X"28",X"02",X"CB",X"DF",X"08",X"21",X"00",X"44",X"CD",X"D2",X"02",X"08",X"CB",
		X"47",X"28",X"02",X"CB",X"E7",X"CB",X"4F",X"28",X"02",X"CB",X"EF",X"08",X"31",X"FD",X"43",X"21",
		X"00",X"4C",X"CD",X"D2",X"02",X"08",X"CB",X"47",X"28",X"02",X"CB",X"F7",X"CB",X"4F",X"28",X"02",
		X"CB",X"FF",X"08",X"3E",X"01",X"CD",X"55",X"15",X"21",X"00",X"40",X"11",X"01",X"40",X"01",X"FE",
		X"03",X"36",X"40",X"ED",X"B0",X"11",X"66",X"41",X"21",X"ED",X"1B",X"3E",X"01",X"06",X"0B",X"CD",
		X"66",X"16",X"11",X"8A",X"40",X"21",X"F8",X"1B",X"3E",X"01",X"06",X"18",X"CD",X"66",X"16",X"11",
		X"EC",X"40",X"21",X"10",X"1C",X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"11",X"ED",X"40",X"21",
		X"24",X"1C",X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"11",X"EE",X"40",X"21",X"38",X"1C",X"3E",
		X"01",X"06",X"14",X"CD",X"66",X"16",X"11",X"EF",X"40",X"21",X"4C",X"1C",X"3E",X"01",X"06",X"14",
		X"CD",X"66",X"16",X"11",X"93",X"40",X"21",X"DC",X"1C",X"3E",X"01",X"06",X"18",X"CD",X"66",X"16",
		X"11",X"F5",X"40",X"21",X"60",X"1C",X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"11",X"F6",X"40",
		X"21",X"74",X"1C",X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"11",X"F7",X"40",X"21",X"88",X"1C",
		X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"11",X"F8",X"40",X"21",X"9C",X"1C",X"3E",X"01",X"06",
		X"14",X"CD",X"66",X"16",X"11",X"F9",X"40",X"21",X"B0",X"1C",X"3E",X"01",X"06",X"14",X"CD",X"66",
		X"16",X"11",X"FA",X"40",X"21",X"C4",X"1C",X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"08",X"32",
		X"FB",X"4D",X"08",X"3A",X"FB",X"4D",X"CB",X"57",X"28",X"0D",X"11",X"F5",X"40",X"21",X"D8",X"1C",
		X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"5F",X"28",X"0D",X"11",X"F6",
		X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"67",
		X"28",X"0D",X"11",X"F7",X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",
		X"FB",X"4D",X"CB",X"6F",X"28",X"0D",X"11",X"F8",X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",
		X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"77",X"28",X"0D",X"11",X"F9",X"40",X"21",X"D8",X"1C",
		X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"7F",X"28",X"0D",X"11",X"FA",
		X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"1E",X"00",X"21",X"00",X"00",
		X"CD",X"B9",X"02",X"30",X"02",X"CB",X"C3",X"21",X"00",X"10",X"CD",X"B9",X"02",X"30",X"02",X"CB",
		X"CB",X"21",X"00",X"20",X"CD",X"B9",X"02",X"30",X"02",X"CB",X"D3",X"21",X"00",X"30",X"CD",X"B9",
		X"02",X"30",X"02",X"CB",X"DB",X"3A",X"FB",X"4D",X"FE",X"00",X"28",X"02",X"3E",X"80",X"B3",X"32",
		X"FB",X"4D",X"CB",X"47",X"28",X"0D",X"11",X"EC",X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",
		X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"4F",X"28",X"0D",X"11",X"ED",X"40",X"21",X"D8",X"1C",
		X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"57",X"28",X"0D",X"11",X"EE",
		X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",X"FB",X"4D",X"CB",X"5F",
		X"28",X"0D",X"11",X"EF",X"40",X"21",X"D8",X"1C",X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"3A",
		X"FB",X"4D",X"FE",X"00",X"20",X"0E",X"FB",X"3E",X"01",X"32",X"00",X"50",X"3E",X"02",X"CD",X"70",
		X"15",X"C3",X"95",X"00",X"32",X"C0",X"50",X"18",X"FB",X"01",X"00",X"10",X"AF",X"32",X"C0",X"50",
		X"86",X"23",X"57",X"0B",X"79",X"B0",X"7A",X"20",X"F7",X"FE",X"FF",X"28",X"02",X"37",X"C9",X"37",
		X"3F",X"C9",X"08",X"E6",X"FC",X"08",X"E5",X"3E",X"11",X"CD",X"F1",X"02",X"E1",X"E5",X"3E",X"22",
		X"CD",X"F1",X"02",X"E1",X"E5",X"3E",X"44",X"CD",X"F1",X"02",X"E1",X"3E",X"88",X"CD",X"F1",X"02",
		X"C9",X"32",X"C0",X"50",X"E5",X"E5",X"D1",X"13",X"01",X"FF",X"03",X"77",X"ED",X"B0",X"E1",X"01",
		X"00",X"04",X"BE",X"C4",X"0F",X"03",X"23",X"5F",X"0B",X"79",X"B0",X"7B",X"20",X"F4",X"C9",X"5F",
		X"7E",X"E6",X"0F",X"57",X"7B",X"E6",X"0F",X"BA",X"28",X"04",X"08",X"CB",X"CF",X"08",X"7E",X"E6",
		X"F0",X"57",X"7B",X"E6",X"F0",X"BA",X"C8",X"08",X"CB",X"C7",X"08",X"7B",X"C9",X"0B",X"4C",X"49",
		X"5A",X"41",X"52",X"44",X"20",X"57",X"49",X"5A",X"41",X"52",X"44",X"2C",X"43",X"4F",X"50",X"59",
		X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"54",X"45",X"43",X"48",X"53",X"54",
		X"41",X"52",X"20",X"49",X"4E",X"43",X"2E",X"32",X"C0",X"50",X"21",X"00",X"40",X"11",X"01",X"40",
		X"01",X"FE",X"07",X"36",X"40",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"00",X"4C",X"11",X"01",X"4C",
		X"01",X"FE",X"03",X"36",X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"60",X"50",X"11",X"61",X"50",
		X"01",X"0F",X"00",X"36",X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"F0",X"4F",X"11",X"F1",X"4F",
		X"01",X"0F",X"00",X"36",X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"40",X"50",X"11",X"41",X"50",
		X"01",X"1F",X"00",X"36",X"00",X"ED",X"B0",X"21",X"A2",X"4C",X"11",X"A3",X"4C",X"01",X"4F",X"00",
		X"36",X"FF",X"ED",X"B0",X"21",X"CB",X"8B",X"22",X"8E",X"4D",X"3A",X"80",X"50",X"47",X"E6",X"03",
		X"32",X"96",X"4D",X"21",X"66",X"1D",X"CD",X"E3",X"15",X"7E",X"32",X"97",X"4D",X"78",X"E6",X"0C",
		X"CB",X"3F",X"CB",X"3F",X"21",X"C7",X"8B",X"CD",X"E3",X"15",X"7E",X"32",X"9D",X"4D",X"78",X"E6",
		X"30",X"21",X"87",X"8B",X"CD",X"E3",X"15",X"22",X"9E",X"4D",X"78",X"E6",X"30",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"32",X"A0",X"4D",X"78",X"CB",X"77",X"20",X"05",X"21",X"91",X"4D",
		X"CB",X"FE",X"ED",X"56",X"FB",X"3E",X"01",X"32",X"00",X"50",X"CD",X"80",X"8A",X"21",X"C2",X"43",
		X"11",X"C3",X"43",X"01",X"3C",X"00",X"36",X"40",X"ED",X"B0",X"21",X"C2",X"47",X"11",X"C3",X"47",
		X"01",X"1C",X"00",X"36",X"1A",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"E2",X"47",X"11",X"E3",X"47",
		X"01",X"1C",X"00",X"36",X"1B",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"9A",X"1A",X"11",X"C3",X"43",
		X"01",X"1A",X"00",X"ED",X"B0",X"AF",X"32",X"E4",X"43",X"32",X"ED",X"43",X"32",X"F6",X"43",X"21",
		X"D4",X"8B",X"11",X"AF",X"4D",X"01",X"3C",X"00",X"ED",X"B0",X"21",X"B4",X"4D",X"11",X"F2",X"43",
		X"CD",X"ED",X"15",X"C3",X"7E",X"04",X"DD",X"7E",X"04",X"80",X"FD",X"96",X"04",X"CB",X"20",X"04",
		X"B8",X"D0",X"DD",X"7E",X"05",X"81",X"FD",X"96",X"05",X"CB",X"21",X"0C",X"B9",X"C9",X"21",X"02",
		X"40",X"11",X"03",X"40",X"01",X"3C",X"00",X"36",X"40",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"02",
		X"44",X"11",X"03",X"44",X"01",X"1C",X"00",X"36",X"01",X"ED",X"B0",X"21",X"02",X"44",X"11",X"03",
		X"44",X"01",X"09",X"00",X"36",X"09",X"ED",X"B0",X"21",X"15",X"44",X"11",X"16",X"44",X"01",X"09",
		X"00",X"36",X"08",X"ED",X"B0",X"21",X"22",X"44",X"11",X"23",X"44",X"01",X"1C",X"00",X"36",X"18",
		X"ED",X"B0",X"32",X"C0",X"50",X"21",X"B4",X"1A",X"11",X"0F",X"40",X"01",X"06",X"00",X"ED",X"B0",
		X"AF",X"32",X"0C",X"40",X"3A",X"96",X"4D",X"FE",X"00",X"20",X"0B",X"21",X"BA",X"1A",X"11",X"0C",
		X"40",X"01",X"09",X"00",X"ED",X"B0",X"32",X"C0",X"50",X"21",X"02",X"4E",X"11",X"03",X"4E",X"01",
		X"F2",X"00",X"36",X"00",X"ED",X"B0",X"21",X"6C",X"8C",X"22",X"1B",X"4E",X"22",X"03",X"4E",X"21",
		X"1A",X"4E",X"22",X"0A",X"4E",X"21",X"9A",X"8C",X"22",X"36",X"4E",X"22",X"1E",X"4E",X"21",X"35",
		X"4E",X"22",X"25",X"4E",X"21",X"B1",X"8C",X"22",X"51",X"4E",X"22",X"39",X"4E",X"21",X"50",X"4E",
		X"22",X"40",X"4E",X"21",X"C9",X"8C",X"22",X"6C",X"4E",X"22",X"54",X"4E",X"21",X"6B",X"4E",X"22",
		X"5B",X"4E",X"21",X"FB",X"8C",X"22",X"87",X"4E",X"22",X"6F",X"4E",X"21",X"86",X"4E",X"22",X"76",
		X"4E",X"21",X"16",X"8D",X"22",X"A2",X"4E",X"22",X"8A",X"4E",X"21",X"A1",X"4E",X"22",X"91",X"4E",
		X"21",X"2C",X"8D",X"22",X"BD",X"4E",X"22",X"A5",X"4E",X"21",X"BC",X"4E",X"22",X"AC",X"4E",X"21",
		X"FC",X"8E",X"22",X"D8",X"4E",X"22",X"C0",X"4E",X"21",X"D7",X"4E",X"22",X"C7",X"4E",X"21",X"14",
		X"8F",X"22",X"F3",X"4E",X"22",X"DB",X"4E",X"21",X"F2",X"4E",X"22",X"E2",X"4E",X"06",X"20",X"21",
		X"40",X"50",X"36",X"00",X"23",X"10",X"FB",X"21",X"91",X"4D",X"CB",X"EE",X"3A",X"96",X"4D",X"FE",
		X"00",X"CA",X"EE",X"06",X"3A",X"95",X"4D",X"FE",X"00",X"C2",X"EE",X"06",X"21",X"90",X"4D",X"CB",
		X"A6",X"AF",X"32",X"01",X"50",X"21",X"91",X"4D",X"CB",X"86",X"CD",X"24",X"12",X"32",X"C0",X"50",
		X"CD",X"69",X"90",X"21",X"90",X"4D",X"CB",X"6E",X"C2",X"EE",X"06",X"CD",X"5D",X"11",X"3E",X"07",
		X"CD",X"70",X"15",X"21",X"90",X"4D",X"CB",X"6E",X"C2",X"EE",X"06",X"3E",X"40",X"CD",X"45",X"15",
		X"11",X"44",X"44",X"21",X"10",X"8C",X"3E",X"01",X"06",X"1C",X"CD",X"7C",X"16",X"11",X"59",X"44",
		X"21",X"12",X"8C",X"3E",X"01",X"06",X"1C",X"CD",X"7C",X"16",X"11",X"5C",X"44",X"21",X"11",X"8C",
		X"3E",X"01",X"06",X"1C",X"CD",X"7C",X"16",X"11",X"44",X"41",X"21",X"83",X"1B",X"3E",X"01",X"06",
		X"0C",X"CD",X"66",X"16",X"CD",X"C9",X"8A",X"3A",X"96",X"4D",X"FE",X"01",X"20",X"0F",X"11",X"19",
		X"41",X"21",X"8F",X"1B",X"3E",X"01",X"06",X"0F",X"CD",X"66",X"16",X"18",X"20",X"FE",X"02",X"20",
		X"0F",X"11",X"19",X"41",X"21",X"9E",X"1B",X"3E",X"01",X"06",X"0F",X"CD",X"66",X"16",X"18",X"0D",
		X"11",X"19",X"41",X"21",X"AD",X"1B",X"3E",X"01",X"06",X"0F",X"CD",X"66",X"16",X"11",X"9C",X"40",
		X"21",X"BC",X"1B",X"3E",X"01",X"06",X"19",X"CD",X"66",X"16",X"3A",X"A0",X"4D",X"FE",X"00",X"20",
		X"0F",X"11",X"7C",X"41",X"21",X"D5",X"1B",X"3E",X"01",X"06",X"06",X"CD",X"66",X"16",X"18",X"33",
		X"FE",X"01",X"20",X"0F",X"11",X"7C",X"41",X"21",X"DB",X"1B",X"3E",X"01",X"06",X"06",X"CD",X"66",
		X"16",X"18",X"20",X"FE",X"02",X"20",X"0F",X"11",X"7C",X"41",X"21",X"E1",X"1B",X"3E",X"01",X"06",
		X"06",X"CD",X"66",X"16",X"18",X"0D",X"11",X"7C",X"41",X"21",X"E7",X"1B",X"3E",X"01",X"06",X"06",
		X"CD",X"66",X"16",X"3E",X"0D",X"CD",X"70",X"15",X"21",X"90",X"4D",X"CB",X"6E",X"20",X"4F",X"CD",
		X"81",X"8A",X"3E",X"0B",X"32",X"FC",X"4D",X"21",X"13",X"8C",X"22",X"FD",X"4D",X"CD",X"9D",X"8A",
		X"21",X"91",X"4D",X"CB",X"EE",X"CD",X"07",X"10",X"CD",X"D2",X"17",X"CD",X"86",X"1D",X"AF",X"32",
		X"1D",X"4E",X"32",X"38",X"4E",X"32",X"53",X"4E",X"32",X"6E",X"4E",X"32",X"89",X"4E",X"32",X"A4",
		X"4E",X"32",X"BF",X"4E",X"32",X"DA",X"4E",X"CD",X"C4",X"15",X"32",X"C0",X"50",X"21",X"90",X"4D",
		X"CB",X"6E",X"20",X"0A",X"21",X"91",X"4D",X"CB",X"6E",X"CA",X"AA",X"05",X"18",X"CA",X"CD",X"24",
		X"12",X"21",X"90",X"4D",X"CB",X"E6",X"CB",X"AE",X"21",X"91",X"4D",X"CB",X"AE",X"CB",X"9E",X"CB",
		X"C6",X"21",X"A2",X"4C",X"11",X"A3",X"4C",X"01",X"4F",X"00",X"36",X"FF",X"ED",X"B0",X"3E",X"FF",
		X"32",X"01",X"50",X"32",X"C0",X"50",X"3E",X"40",X"CD",X"45",X"15",X"3E",X"1B",X"CD",X"55",X"15",
		X"3A",X"96",X"4D",X"FE",X"00",X"CA",X"B4",X"07",X"3A",X"95",X"4D",X"FE",X"02",X"30",X"55",X"11",
		X"78",X"41",X"21",X"C3",X"1A",X"3E",X"01",X"06",X"0B",X"CD",X"66",X"16",X"CD",X"C9",X"8A",X"3A",
		X"40",X"50",X"CB",X"6F",X"C2",X"C7",X"07",X"3A",X"96",X"4D",X"FE",X"00",X"28",X"15",X"3A",X"95",
		X"4D",X"FE",X"02",X"38",X"72",X"D6",X"02",X"32",X"95",X"4D",X"3A",X"98",X"4D",X"D6",X"01",X"27",
		X"32",X"98",X"4D",X"21",X"91",X"4D",X"CB",X"E6",X"3A",X"9D",X"4D",X"32",X"A1",X"4D",X"CD",X"06",
		X"00",X"21",X"91",X"4D",X"CB",X"EE",X"3A",X"96",X"4D",X"FE",X"00",X"CA",X"0F",X"08",X"CD",X"36",
		X"11",X"C3",X"0F",X"08",X"FE",X"04",X"30",X"2C",X"11",X"18",X"41",X"21",X"CE",X"1A",X"3E",X"01",
		X"06",X"11",X"CD",X"66",X"16",X"11",X"1A",X"42",X"21",X"DF",X"1A",X"3E",X"01",X"06",X"02",X"CD",
		X"66",X"16",X"11",X"7C",X"41",X"21",X"C3",X"1A",X"3E",X"01",X"06",X"0B",X"CD",X"66",X"16",X"CD",
		X"C9",X"8A",X"18",X"8B",X"11",X"9A",X"40",X"21",X"E1",X"1A",X"3E",X"01",X"06",X"19",X"CD",X"66",
		X"16",X"CD",X"C9",X"8A",X"C3",X"3F",X"07",X"3A",X"40",X"50",X"CB",X"77",X"20",X"2F",X"3A",X"96",
		X"4D",X"FE",X"00",X"28",X"15",X"3A",X"95",X"4D",X"FE",X"04",X"38",X"21",X"D6",X"04",X"32",X"95",
		X"4D",X"3A",X"98",X"4D",X"D6",X"02",X"27",X"32",X"98",X"4D",X"21",X"91",X"4D",X"CB",X"A6",X"3A",
		X"9D",X"4D",X"32",X"A2",X"4D",X"CB",X"CE",X"CD",X"3B",X"00",X"C3",X"68",X"07",X"32",X"C0",X"50",
		X"21",X"90",X"4D",X"CB",X"76",X"20",X"03",X"C3",X"3F",X"07",X"CB",X"B6",X"C3",X"13",X"07",X"AF",
		X"21",X"A3",X"4D",X"11",X"A4",X"4D",X"01",X"09",X"00",X"77",X"ED",X"B0",X"32",X"AD",X"4D",X"32",
		X"AE",X"4D",X"3E",X"40",X"21",X"E4",X"43",X"11",X"E5",X"43",X"01",X"05",X"00",X"77",X"ED",X"B0",
		X"21",X"F6",X"43",X"11",X"F7",X"43",X"01",X"05",X"00",X"77",X"ED",X"B0",X"AF",X"32",X"E4",X"43",
		X"32",X"F6",X"43",X"AF",X"32",X"FC",X"4D",X"CD",X"A3",X"8A",X"21",X"DA",X"4E",X"CB",X"C6",X"21",
		X"91",X"4D",X"CB",X"66",X"20",X"0A",X"3A",X"A2",X"4D",X"3D",X"32",X"A2",X"4D",X"CD",X"3B",X"00",
		X"3A",X"A1",X"4D",X"3D",X"32",X"A1",X"4D",X"CD",X"06",X"00",X"CD",X"07",X"10",X"CD",X"57",X"85",
		X"32",X"C0",X"50",X"3A",X"DA",X"4E",X"FE",X"00",X"20",X"F6",X"CD",X"86",X"1D",X"21",X"92",X"4D",
		X"CB",X"66",X"28",X"13",X"CB",X"A6",X"ED",X"5B",X"A9",X"4D",X"7B",X"B2",X"28",X"1C",X"21",X"00",
		X"00",X"22",X"A9",X"4D",X"C3",X"A7",X"08",X"CB",X"E6",X"ED",X"5B",X"AB",X"4D",X"7B",X"B2",X"28",
		X"09",X"21",X"00",X"00",X"22",X"AB",X"4D",X"CD",X"7A",X"10",X"32",X"C0",X"50",X"CD",X"C4",X"15",
		X"21",X"91",X"4D",X"CB",X"6E",X"C2",X"D6",X"09",X"CB",X"4E",X"C2",X"D6",X"09",X"CD",X"CD",X"89",
		X"CD",X"24",X"12",X"ED",X"5B",X"A9",X"4D",X"7B",X"B2",X"28",X"0E",X"21",X"00",X"00",X"22",X"A9",
		X"4D",X"21",X"92",X"4D",X"CB",X"A6",X"CD",X"7A",X"10",X"ED",X"5B",X"AB",X"4D",X"7B",X"B2",X"28",
		X"0E",X"21",X"00",X"00",X"22",X"AB",X"4D",X"21",X"92",X"4D",X"CB",X"E6",X"CD",X"7A",X"10",X"DD",
		X"21",X"00",X"4E",X"21",X"91",X"4D",X"CB",X"6E",X"20",X"0A",X"3A",X"A1",X"4D",X"B7",X"20",X"04",
		X"DD",X"CB",X"00",X"C6",X"CB",X"4E",X"20",X"0E",X"CB",X"66",X"20",X"0A",X"3A",X"A2",X"4D",X"B7",
		X"20",X"04",X"DD",X"CB",X"00",X"CE",X"DD",X"7E",X"00",X"B7",X"28",X"69",X"CD",X"65",X"15",X"11",
		X"6F",X"41",X"21",X"C3",X"1A",X"3E",X"01",X"06",X"0B",X"CD",X"66",X"16",X"11",X"31",X"41",X"21",
		X"F4",X"1C",X"3E",X"01",X"06",X"0F",X"CD",X"66",X"16",X"DD",X"7E",X"00",X"FE",X"03",X"28",X"20",
		X"CB",X"47",X"28",X"0F",X"11",X"6D",X"41",X"21",X"FD",X"1A",X"3E",X"01",X"06",X"0A",X"CD",X"66",
		X"16",X"18",X"0D",X"11",X"6D",X"41",X"21",X"0A",X"1B",X"3E",X"01",X"06",X"0A",X"CD",X"66",X"16",
		X"3E",X"02",X"CD",X"CE",X"15",X"DD",X"7E",X"01",X"3C",X"DD",X"77",X"01",X"FE",X"96",X"20",X"0D",
		X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",X"CD",X"65",X"15",X"18",X"08",X"DD",X"7E",X"00",
		X"B7",X"20",X"DD",X"18",X"EB",X"21",X"91",X"4D",X"CB",X"6E",X"20",X"13",X"3A",X"A1",X"4D",X"FE",
		X"00",X"28",X"0C",X"3D",X"32",X"A1",X"4D",X"CD",X"06",X"00",X"21",X"91",X"4D",X"CB",X"EE",X"CB",
		X"4E",X"20",X"13",X"3A",X"A2",X"4D",X"FE",X"00",X"28",X"34",X"3D",X"32",X"A2",X"4D",X"CD",X"3B",
		X"00",X"21",X"91",X"4D",X"CB",X"CE",X"CB",X"5E",X"CA",X"6A",X"08",X"CB",X"9E",X"21",X"92",X"4D",
		X"CB",X"CE",X"3A",X"FC",X"4D",X"FE",X"0F",X"28",X"04",X"3C",X"32",X"FC",X"4D",X"CD",X"CE",X"89",
		X"CD",X"CC",X"89",X"C3",X"6A",X"08",X"CB",X"5E",X"C2",X"BD",X"08",X"C3",X"7A",X"08",X"CB",X"6E",
		X"C2",X"B6",X"09",X"CD",X"65",X"15",X"11",X"90",X"41",X"21",X"14",X"1B",X"3E",X"01",X"06",X"09",
		X"CD",X"66",X"16",X"3E",X"02",X"CD",X"70",X"15",X"CD",X"38",X"12",X"21",X"90",X"4D",X"CB",X"F6",
		X"21",X"91",X"4D",X"CB",X"9E",X"C3",X"87",X"05",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"AF",X"32",X"00",X"50",X"2A",X"8E",X"4D",X"23",X"22",X"8E",X"4D",X"7E",X"FE",X"FF",X"C2",X"27",
		X"0A",X"21",X"CB",X"8B",X"22",X"8E",X"4D",X"2A",X"A2",X"4C",X"3A",X"A4",X"4C",X"77",X"2A",X"A5",
		X"4C",X"3A",X"A7",X"4C",X"77",X"2A",X"AA",X"4C",X"3A",X"AC",X"4C",X"77",X"2A",X"AD",X"4C",X"3A",
		X"AF",X"4C",X"77",X"2A",X"B2",X"4C",X"3A",X"B4",X"4C",X"77",X"2A",X"B5",X"4C",X"3A",X"B7",X"4C",
		X"77",X"2A",X"BA",X"4C",X"3A",X"BC",X"4C",X"77",X"2A",X"BD",X"4C",X"3A",X"BF",X"4C",X"77",X"2A",
		X"C2",X"4C",X"3A",X"C4",X"4C",X"77",X"2A",X"C5",X"4C",X"3A",X"C7",X"4C",X"77",X"2A",X"CA",X"4C",
		X"3A",X"CC",X"4C",X"77",X"2A",X"CD",X"4C",X"3A",X"CF",X"4C",X"77",X"2A",X"D2",X"4C",X"3A",X"D4",
		X"4C",X"77",X"2A",X"D5",X"4C",X"3A",X"D7",X"4C",X"77",X"2A",X"DA",X"4C",X"3A",X"DC",X"4C",X"77",
		X"2A",X"DD",X"4C",X"3A",X"DF",X"4C",X"77",X"2A",X"E2",X"4C",X"3A",X"E4",X"4C",X"77",X"2A",X"E5",
		X"4C",X"3A",X"E7",X"4C",X"77",X"2A",X"EA",X"4C",X"3A",X"EC",X"4C",X"77",X"2A",X"ED",X"4C",X"3A",
		X"EF",X"4C",X"77",X"ED",X"5B",X"FD",X"4C",X"CD",X"F8",X"0D",X"ED",X"53",X"62",X"50",X"ED",X"5B",
		X"15",X"4D",X"CD",X"F8",X"0D",X"ED",X"53",X"64",X"50",X"ED",X"5B",X"2D",X"4D",X"CD",X"F8",X"0D",
		X"ED",X"53",X"66",X"50",X"ED",X"5B",X"45",X"4D",X"CD",X"F8",X"0D",X"ED",X"53",X"68",X"50",X"ED",
		X"5B",X"5D",X"4D",X"CD",X"F8",X"0D",X"ED",X"53",X"6A",X"50",X"ED",X"5B",X"75",X"4D",X"CD",X"F8",
		X"0D",X"ED",X"53",X"6C",X"50",X"2A",X"FF",X"4C",X"CD",X"11",X"0E",X"22",X"F2",X"4F",X"2A",X"17",
		X"4D",X"CD",X"11",X"0E",X"22",X"F4",X"4F",X"2A",X"2F",X"4D",X"CD",X"11",X"0E",X"22",X"F6",X"4F",
		X"2A",X"47",X"4D",X"CD",X"11",X"0E",X"22",X"F8",X"4F",X"2A",X"5F",X"4D",X"CD",X"11",X"0E",X"22",
		X"FA",X"4F",X"2A",X"77",X"4D",X"CD",X"11",X"0E",X"22",X"FC",X"4F",X"21",X"90",X"4D",X"CB",X"46",
		X"20",X"58",X"3A",X"00",X"50",X"CB",X"6F",X"CA",X"FB",X"0B",X"CB",X"8E",X"CB",X"56",X"20",X"3F",
		X"3A",X"00",X"50",X"CB",X"7F",X"CA",X"09",X"0C",X"3A",X"93",X"4D",X"FE",X"06",X"28",X"07",X"3C",
		X"32",X"93",X"4D",X"C3",X"0E",X"0C",X"AF",X"32",X"93",X"4D",X"CB",X"5E",X"20",X"0A",X"3A",X"94",
		X"4D",X"FE",X"00",X"20",X"0C",X"C3",X"0E",X"0C",X"AF",X"32",X"07",X"50",X"CB",X"9E",X"C3",X"0E",
		X"0C",X"3D",X"32",X"94",X"4D",X"3E",X"01",X"32",X"07",X"50",X"CB",X"DE",X"C3",X"0E",X"0C",X"3A",
		X"00",X"50",X"CB",X"7F",X"28",X"C2",X"CB",X"96",X"18",X"10",X"3A",X"00",X"50",X"CB",X"6F",X"28",
		X"AB",X"CB",X"86",X"3A",X"94",X"4D",X"3C",X"32",X"94",X"4D",X"3A",X"00",X"4E",X"B7",X"28",X"2A",
		X"CB",X"47",X"28",X"0D",X"CB",X"87",X"32",X"00",X"4E",X"3E",X"02",X"32",X"A1",X"4D",X"CD",X"06",
		X"00",X"3A",X"00",X"4E",X"CB",X"4F",X"28",X"36",X"CB",X"8F",X"32",X"00",X"4E",X"3E",X"02",X"32",
		X"A2",X"4D",X"CD",X"3B",X"00",X"21",X"90",X"4D",X"18",X"24",X"21",X"90",X"4D",X"3A",X"95",X"4D",
		X"FE",X"14",X"30",X"1A",X"47",X"3A",X"97",X"4D",X"80",X"32",X"95",X"4D",X"CB",X"3F",X"06",X"00",
		X"80",X"27",X"32",X"98",X"4D",X"CD",X"36",X"11",X"CB",X"66",X"20",X"02",X"CB",X"EE",X"3A",X"02",
		X"4E",X"CB",X"C7",X"32",X"02",X"4E",X"CB",X"F6",X"C3",X"48",X"0B",X"CB",X"4E",X"20",X"05",X"CB",
		X"CE",X"C3",X"3C",X"0B",X"CB",X"C6",X"C3",X"3A",X"0B",X"CB",X"D6",X"C3",X"48",X"0B",X"00",X"21",
		X"91",X"4D",X"CB",X"46",X"28",X"09",X"CD",X"35",X"18",X"CD",X"15",X"18",X"CD",X"25",X"18",X"3A",
		X"9A",X"4D",X"3C",X"32",X"9A",X"4D",X"3A",X"99",X"4D",X"3C",X"32",X"99",X"4D",X"FE",X"3C",X"20",
		X"0B",X"AF",X"32",X"99",X"4D",X"3A",X"9B",X"4D",X"3C",X"32",X"9B",X"4D",X"21",X"90",X"4D",X"CB",
		X"BE",X"3A",X"00",X"50",X"CB",X"77",X"20",X"35",X"AF",X"32",X"01",X"50",X"21",X"62",X"50",X"06",
		X"0C",X"36",X"00",X"23",X"10",X"FB",X"3E",X"40",X"CD",X"45",X"15",X"3E",X"02",X"CD",X"55",X"15",
		X"11",X"D0",X"41",X"21",X"7F",X"1B",X"3E",X"01",X"06",X"04",X"CD",X"66",X"16",X"06",X"FF",X"21",
		X"FF",X"FF",X"2B",X"7D",X"BC",X"32",X"C0",X"50",X"20",X"F8",X"10",X"F3",X"76",X"FB",X"3E",X"01",
		X"32",X"00",X"50",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"ED",X"4D",X"DD",X"2A",X"89",
		X"4D",X"DD",X"7E",X"00",X"CB",X"27",X"21",X"E4",X"0C",X"CD",X"E3",X"15",X"23",X"7E",X"32",X"8B",
		X"4D",X"2B",X"DD",X"7E",X"03",X"32",X"8C",X"4D",X"DD",X"7E",X"05",X"32",X"8D",X"4D",X"7E",X"FE",
		X"00",X"28",X"0F",X"CD",X"24",X"0D",X"3A",X"8C",X"4D",X"DD",X"77",X"03",X"3A",X"8D",X"4D",X"DD",
		X"77",X"05",X"DD",X"7E",X"02",X"32",X"8C",X"4D",X"DD",X"7E",X"04",X"32",X"8D",X"4D",X"3A",X"8B",
		X"4D",X"FE",X"00",X"C8",X"CD",X"24",X"0D",X"3A",X"8C",X"4D",X"DD",X"77",X"02",X"3A",X"8D",X"4D",
		X"DD",X"77",X"04",X"C9",X"04",X"00",X"04",X"06",X"04",X"0A",X"04",X"0E",X"04",X"02",X"10",X"02",
		X"0C",X"02",X"08",X"02",X"00",X"02",X"06",X"02",X"0A",X"02",X"0E",X"02",X"02",X"02",X"02",X"0E",
		X"02",X"0A",X"02",X"06",X"02",X"00",X"02",X"08",X"02",X"0C",X"02",X"10",X"02",X"04",X"0E",X"04",
		X"0A",X"04",X"06",X"04",X"00",X"04",X"08",X"04",X"0C",X"04",X"10",X"04",X"04",X"04",X"04",X"10",
		X"04",X"0C",X"04",X"08",X"11",X"44",X"0D",X"CD",X"E8",X"15",X"1A",X"6F",X"13",X"1A",X"67",X"E9",
		X"3A",X"8C",X"4D",X"80",X"47",X"E6",X"0F",X"32",X"8C",X"4D",X"CB",X"38",X"CB",X"38",X"CB",X"38",
		X"CB",X"38",X"3A",X"8D",X"4D",X"C9",X"56",X"0D",X"61",X"0D",X"6C",X"0D",X"7B",X"0D",X"8A",X"0D",
		X"97",X"0D",X"A4",X"0D",X"BA",X"0D",X"DD",X"46",X"01",X"CD",X"30",X"0D",X"80",X"32",X"8D",X"4D",
		X"C9",X"DD",X"46",X"01",X"CD",X"30",X"0D",X"90",X"32",X"8D",X"4D",X"C9",X"DD",X"46",X"01",X"CB",
		X"38",X"CB",X"38",X"CD",X"30",X"0D",X"80",X"32",X"8D",X"4D",X"C9",X"DD",X"46",X"01",X"CB",X"38",
		X"CB",X"38",X"CD",X"30",X"0D",X"90",X"32",X"8D",X"4D",X"C9",X"DD",X"46",X"01",X"CB",X"38",X"CD",
		X"30",X"0D",X"80",X"32",X"8D",X"4D",X"C9",X"DD",X"46",X"01",X"CB",X"38",X"CD",X"30",X"0D",X"90",
		X"32",X"8D",X"4D",X"C9",X"DD",X"46",X"01",X"CB",X"38",X"CB",X"38",X"DD",X"7E",X"01",X"CB",X"3F",
		X"80",X"47",X"CD",X"30",X"0D",X"80",X"32",X"8D",X"4D",X"C9",X"DD",X"46",X"01",X"CB",X"38",X"CB",
		X"38",X"DD",X"7E",X"01",X"CB",X"3F",X"80",X"47",X"CD",X"30",X"0D",X"90",X"32",X"8D",X"4D",X"C9",
		X"3A",X"F2",X"4C",X"E6",X"07",X"32",X"A0",X"4C",X"3A",X"F3",X"4C",X"E6",X"07",X"32",X"A1",X"4C",
		X"3A",X"F2",X"4C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"57",X"3A",X"F3",X"4C",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"5F",X"CD",X"58",X"10",X"C9",X"D5",X"37",X"3F",X"21",X"0E",X"01",X"16",X"00",
		X"ED",X"52",X"7D",X"37",X"3F",X"21",X"10",X"01",X"D1",X"5A",X"16",X"00",X"ED",X"52",X"55",X"5F",
		X"C9",X"7D",X"EE",X"03",X"6F",X"C9",X"2A",X"F4",X"4C",X"EB",X"DD",X"21",X"00",X"00",X"DD",X"19",
		X"EB",X"01",X"00",X"4C",X"37",X"3F",X"ED",X"42",X"CB",X"3C",X"CB",X"1D",X"E5",X"DD",X"7E",X"00",
		X"21",X"3D",X"0E",X"CB",X"27",X"CD",X"E3",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"0F",X"0F",X"49",
		X"0E",X"8E",X"0E",X"1E",X"0F",X"28",X"0F",X"3B",X"0F",X"F3",X"DD",X"7E",X"04",X"32",X"F2",X"4C",
		X"DD",X"7E",X"03",X"32",X"F3",X"4C",X"CD",X"D0",X"0D",X"DD",X"7E",X"06",X"12",X"3A",X"A0",X"4C",
		X"FE",X"00",X"20",X"18",X"3A",X"A1",X"4C",X"FE",X"00",X"20",X"18",X"C1",X"21",X"A2",X"4C",X"09",
		X"E5",X"D1",X"13",X"01",X"05",X"00",X"36",X"FF",X"ED",X"B0",X"FB",X"C9",X"DD",X"7E",X"06",X"13",
		X"12",X"18",X"E8",X"DD",X"7E",X"06",X"21",X"20",X"00",X"19",X"EB",X"12",X"18",X"DD",X"CD",X"B2",
		X"0F",X"DD",X"7E",X"04",X"90",X"32",X"F2",X"4C",X"DD",X"7E",X"03",X"32",X"F3",X"4C",X"CD",X"D0",
		X"0D",X"3A",X"A0",X"4C",X"FE",X"00",X"28",X"32",X"3A",X"A0",X"4C",X"CB",X"27",X"DD",X"46",X"05",
		X"80",X"3D",X"C1",X"FD",X"21",X"A2",X"4C",X"FD",X"09",X"FD",X"73",X"00",X"FD",X"72",X"01",X"FD",
		X"77",X"02",X"3C",X"13",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"77",X"05",X"3A",X"F2",X"4C",
		X"DD",X"77",X"04",X"3A",X"F3",X"4C",X"DD",X"77",X"03",X"C9",X"3A",X"A1",X"4C",X"FE",X"00",X"CA",
		X"44",X"0F",X"3A",X"A1",X"4C",X"CB",X"27",X"C6",X"0F",X"DD",X"46",X"05",X"80",X"C1",X"FD",X"21",
		X"A2",X"4C",X"FD",X"09",X"FD",X"73",X"00",X"FD",X"72",X"01",X"FD",X"77",X"02",X"3C",X"21",X"20",
		X"00",X"19",X"EB",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"77",X"05",X"C3",X"CD",X"0E",X"DD",
		X"7E",X"04",X"32",X"F2",X"4C",X"DD",X"7E",X"03",X"32",X"F3",X"4C",X"C3",X"9E",X"0E",X"CD",X"B2",
		X"0F",X"DD",X"7E",X"04",X"80",X"C3",X"95",X"0E",X"CD",X"B2",X"0F",X"DD",X"7E",X"03",X"90",X"32",
		X"F3",X"4C",X"DD",X"7E",X"04",X"32",X"F2",X"4C",X"C3",X"9E",X"0E",X"CD",X"B2",X"0F",X"DD",X"7E",
		X"03",X"80",X"18",X"EB",X"DD",X"7E",X"05",X"C1",X"FD",X"21",X"A2",X"4C",X"FD",X"09",X"FD",X"73",
		X"00",X"FD",X"72",X"01",X"FD",X"77",X"02",X"3A",X"F2",X"4C",X"DD",X"77",X"04",X"3A",X"F3",X"4C",
		X"DD",X"77",X"03",X"DD",X"7E",X"00",X"21",X"78",X"0F",X"CB",X"27",X"CD",X"E3",X"15",X"D5",X"5E",
		X"23",X"56",X"EB",X"D1",X"DD",X"7E",X"06",X"E9",X"A5",X"0F",X"84",X"0F",X"85",X"0F",X"90",X"0F",
		X"93",X"0F",X"9A",X"0F",X"C9",X"13",X"FD",X"73",X"03",X"FD",X"72",X"04",X"FD",X"77",X"05",X"C9",
		X"1B",X"18",X"F3",X"21",X"20",X"00",X"19",X"EB",X"18",X"EC",X"EB",X"11",X"20",X"00",X"37",X"3F",
		X"ED",X"52",X"EB",X"18",X"E1",X"FD",X"36",X"03",X"FF",X"FD",X"36",X"04",X"FF",X"FD",X"36",X"05",
		X"FF",X"C9",X"DD",X"7E",X"01",X"DD",X"86",X"02",X"47",X"E6",X"0F",X"DD",X"77",X"02",X"CB",X"38",
		X"CB",X"38",X"CB",X"38",X"CB",X"38",X"C9",X"21",X"AF",X"4D",X"11",X"6A",X"42",X"CD",X"78",X"00",
		X"11",X"6C",X"42",X"CD",X"78",X"00",X"11",X"6E",X"42",X"CD",X"78",X"00",X"11",X"70",X"42",X"CD",
		X"78",X"00",X"11",X"72",X"42",X"CD",X"78",X"00",X"11",X"74",X"42",X"CD",X"78",X"00",X"11",X"76",
		X"42",X"CD",X"78",X"00",X"11",X"78",X"42",X"CD",X"78",X"00",X"11",X"7A",X"42",X"CD",X"78",X"00",
		X"11",X"7C",X"42",X"CD",X"78",X"00",X"C9",X"CD",X"00",X"80",X"3A",X"FC",X"4D",X"21",X"18",X"10",
		X"CB",X"27",X"CB",X"27",X"CD",X"E3",X"15",X"E9",X"CD",X"5A",X"81",X"C9",X"CD",X"96",X"81",X"C9",
		X"CD",X"CB",X"81",X"C9",X"CD",X"05",X"82",X"C9",X"CD",X"A1",X"82",X"C9",X"CD",X"78",X"83",X"C9",
		X"CD",X"B2",X"83",X"C9",X"CD",X"E4",X"83",X"C9",X"CD",X"1A",X"84",X"C9",X"CD",X"40",X"84",X"C9",
		X"CD",X"55",X"84",X"C9",X"CD",X"88",X"84",X"C9",X"CD",X"C9",X"84",X"C9",X"CD",X"F1",X"84",X"C9",
		X"CD",X"24",X"85",X"C9",X"CD",X"40",X"85",X"C9",X"D5",X"AF",X"CB",X"23",X"17",X"CB",X"23",X"17",
		X"CB",X"23",X"17",X"CB",X"23",X"17",X"CB",X"23",X"17",X"57",X"EB",X"01",X"40",X"40",X"09",X"06",
		X"00",X"D1",X"4A",X"09",X"EB",X"ED",X"53",X"F6",X"4C",X"C9",X"21",X"91",X"4D",X"CB",X"46",X"C8",
		X"21",X"92",X"4D",X"CB",X"66",X"20",X"43",X"21",X"A3",X"4D",X"7B",X"86",X"27",X"77",X"23",X"7A",
		X"8E",X"27",X"77",X"23",X"3E",X"00",X"8E",X"27",X"77",X"38",X"02",X"18",X"32",X"21",X"92",X"4D",
		X"CB",X"66",X"20",X"13",X"21",X"F6",X"43",X"11",X"F7",X"43",X"01",X"05",X"00",X"36",X"40",X"ED",
		X"B0",X"AF",X"32",X"F6",X"43",X"18",X"18",X"21",X"E4",X"43",X"11",X"E5",X"43",X"01",X"05",X"00",
		X"36",X"40",X"ED",X"B0",X"AF",X"32",X"E4",X"43",X"18",X"05",X"21",X"A6",X"4D",X"18",X"BB",X"21",
		X"92",X"4D",X"CB",X"66",X"20",X"55",X"21",X"A5",X"4D",X"11",X"FB",X"43",X"3A",X"AD",X"4D",X"F5",
		X"CD",X"ED",X"15",X"23",X"23",X"23",X"EB",X"2A",X"9E",X"4D",X"F1",X"FE",X"04",X"D0",X"CB",X"27",
		X"CB",X"27",X"3C",X"3C",X"CD",X"E3",X"15",X"CD",X"03",X"1D",X"D0",X"21",X"1D",X"4E",X"CB",X"C6",
		X"21",X"92",X"4D",X"CB",X"66",X"20",X"12",X"3A",X"AD",X"4D",X"3C",X"32",X"AD",X"4D",X"3A",X"A1",
		X"4D",X"3C",X"32",X"A1",X"4D",X"CD",X"06",X"00",X"C9",X"3A",X"AE",X"4D",X"3C",X"32",X"AE",X"4D",
		X"3A",X"A2",X"4D",X"3C",X"32",X"A2",X"4D",X"CD",X"3B",X"00",X"C9",X"21",X"A8",X"4D",X"11",X"E9",
		X"43",X"3A",X"AE",X"4D",X"18",X"A9",X"3A",X"96",X"4D",X"FE",X"00",X"C8",X"3A",X"98",X"4D",X"E6",
		X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FE",X"00",X"28",X"0C",X"32",X"0D",X"40",
		X"3A",X"98",X"4D",X"E6",X"0F",X"32",X"0C",X"40",X"C9",X"3E",X"40",X"18",X"F0",X"3E",X"40",X"CD",
		X"45",X"15",X"3E",X"02",X"CD",X"55",X"15",X"11",X"29",X"45",X"21",X"9B",X"11",X"3E",X"15",X"06",
		X"0B",X"CD",X"7C",X"16",X"11",X"05",X"41",X"21",X"1D",X"1B",X"3E",X"01",X"06",X"10",X"CD",X"66",
		X"16",X"21",X"29",X"1D",X"11",X"CA",X"42",X"01",X"FF",X"09",X"ED",X"A0",X"13",X"10",X"FB",X"AF",
		X"12",X"CD",X"88",X"15",X"3E",X"01",X"12",X"CD",X"C7",X"0F",X"C9",X"18",X"3E",X"03",X"F5",X"7E",
		X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"3A",X"91",X"4D",X"CB",X"77",
		X"28",X"2A",X"78",X"12",X"3E",X"20",X"CD",X"52",X"16",X"7E",X"E6",X"0F",X"47",X"3A",X"91",X"4D",
		X"CB",X"77",X"32",X"91",X"4D",X"28",X"24",X"78",X"12",X"2B",X"3E",X"20",X"CD",X"52",X"16",X"F1",
		X"3D",X"20",X"CB",X"3A",X"91",X"4D",X"CB",X"B7",X"32",X"91",X"4D",X"C9",X"78",X"FE",X"00",X"28",
		X"D3",X"3A",X"91",X"4D",X"CB",X"F7",X"32",X"91",X"4D",X"18",X"C7",X"78",X"FE",X"00",X"28",X"D9",
		X"3A",X"91",X"4D",X"CB",X"F7",X"32",X"91",X"4D",X"18",X"CD",X"05",X"4C",X"49",X"5A",X"41",X"52",
		X"44",X"20",X"57",X"49",X"5A",X"41",X"52",X"44",X"2C",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",
		X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"54",X"45",X"43",X"48",X"53",X"54",X"41",X"52",X"20",
		X"49",X"4E",X"43",X"2E",X"21",X"F9",X"4C",X"11",X"10",X"00",X"3E",X"06",X"06",X"08",X"36",X"00",
		X"23",X"10",X"FB",X"3D",X"C8",X"19",X"18",X"F4",X"21",X"92",X"4D",X"CB",X"A6",X"21",X"A3",X"4D",
		X"11",X"F1",X"4D",X"01",X"03",X"00",X"ED",X"B0",X"3A",X"F5",X"4D",X"32",X"F4",X"4D",X"CD",X"71",
		X"12",X"21",X"91",X"4D",X"CB",X"66",X"C0",X"21",X"92",X"4D",X"CB",X"E6",X"21",X"A6",X"4D",X"11",
		X"F1",X"4D",X"01",X"03",X"00",X"ED",X"B0",X"3A",X"F6",X"4D",X"32",X"F4",X"4D",X"CD",X"71",X"12",
		X"C9",X"01",X"00",X"0A",X"21",X"ED",X"4D",X"11",X"F3",X"4D",X"2B",X"2B",X"2B",X"C5",X"CD",X"03",
		X"1D",X"C1",X"30",X"0A",X"3E",X"06",X"81",X"4F",X"10",X"ED",X"2B",X"2B",X"18",X"08",X"79",X"FE",
		X"00",X"C8",X"23",X"23",X"23",X"23",X"C5",X"E5",X"06",X"00",X"21",X"EA",X"4D",X"11",X"F0",X"4D",
		X"ED",X"B8",X"3E",X"40",X"CD",X"45",X"15",X"21",X"92",X"4D",X"CB",X"66",X"28",X"0F",X"11",X"62",
		X"41",X"21",X"0A",X"1B",X"3E",X"01",X"06",X"0A",X"CD",X"66",X"16",X"18",X"0D",X"11",X"62",X"41",
		X"21",X"FD",X"1A",X"3E",X"01",X"06",X"0A",X"CD",X"66",X"16",X"11",X"40",X"44",X"21",X"41",X"15",
		X"3E",X"0B",X"06",X"1C",X"CD",X"7C",X"16",X"11",X"4C",X"44",X"21",X"42",X"15",X"3E",X"03",X"06",
		X"1C",X"CD",X"7C",X"16",X"11",X"51",X"44",X"21",X"43",X"15",X"3E",X"10",X"06",X"1C",X"CD",X"7C",
		X"16",X"11",X"50",X"44",X"21",X"44",X"15",X"3E",X"02",X"06",X"1C",X"CD",X"7C",X"16",X"D1",X"D5",
		X"3E",X"40",X"D5",X"E1",X"13",X"01",X"03",X"00",X"77",X"ED",X"B0",X"36",X"00",X"01",X"02",X"00",
		X"ED",X"B0",X"D1",X"C1",X"D5",X"78",X"21",X"6A",X"1D",X"CB",X"27",X"CD",X"E3",X"15",X"4E",X"23",
		X"46",X"C5",X"21",X"80",X"04",X"09",X"0E",X"1A",X"06",X"0F",X"71",X"3E",X"20",X"CD",X"48",X"16",
		X"10",X"F8",X"11",X"C3",X"40",X"21",X"2D",X"1B",X"3E",X"01",X"06",X"14",X"CD",X"66",X"16",X"11",
		X"A5",X"41",X"21",X"41",X"1B",X"3E",X"01",X"06",X"07",X"CD",X"66",X"16",X"11",X"A7",X"40",X"21",
		X"48",X"1B",X"3E",X"01",X"06",X"16",X"CD",X"66",X"16",X"11",X"A8",X"40",X"21",X"5E",X"1B",X"3E",
		X"01",X"06",X"16",X"CD",X"66",X"16",X"11",X"69",X"42",X"21",X"74",X"1B",X"3E",X"01",X"06",X"08",
		X"CD",X"66",X"16",X"11",X"4C",X"40",X"21",X"7C",X"1B",X"3E",X"03",X"06",X"01",X"CD",X"66",X"16",
		X"11",X"8D",X"40",X"21",X"4C",X"1D",X"3E",X"01",X"06",X"1A",X"CD",X"66",X"16",X"3E",X"1A",X"11",
		X"AD",X"47",X"12",X"AF",X"32",X"F7",X"4D",X"32",X"F8",X"4D",X"21",X"AD",X"47",X"22",X"F9",X"4D",
		X"11",X"31",X"41",X"21",X"1D",X"1B",X"3E",X"01",X"06",X"10",X"CD",X"66",X"16",X"21",X"29",X"1D",
		X"11",X"F4",X"42",X"01",X"09",X"00",X"ED",X"B0",X"AF",X"12",X"CD",X"88",X"15",X"3E",X"01",X"12",
		X"21",X"AF",X"4D",X"11",X"94",X"42",X"CD",X"78",X"00",X"11",X"95",X"42",X"CD",X"78",X"00",X"11",
		X"96",X"42",X"CD",X"78",X"00",X"11",X"97",X"42",X"CD",X"78",X"00",X"11",X"98",X"42",X"CD",X"78",
		X"00",X"11",X"99",X"42",X"CD",X"78",X"00",X"11",X"9A",X"42",X"CD",X"78",X"00",X"11",X"9B",X"42",
		X"CD",X"78",X"00",X"11",X"9C",X"42",X"CD",X"78",X"00",X"11",X"9D",X"42",X"CD",X"78",X"00",X"3A",
		X"F5",X"4D",X"21",X"92",X"4D",X"CB",X"66",X"28",X"03",X"3A",X"F6",X"4D",X"CB",X"4F",X"CA",X"9F",
		X"14",X"CB",X"57",X"CA",X"D7",X"14",X"3A",X"F5",X"4D",X"21",X"92",X"4D",X"CB",X"66",X"28",X"03",
		X"3A",X"F6",X"4D",X"CB",X"67",X"C2",X"18",X"15",X"3A",X"F7",X"4D",X"FE",X"1B",X"28",X"1F",X"21",
		X"32",X"1D",X"CD",X"E3",X"15",X"7E",X"E1",X"D1",X"12",X"13",X"77",X"3E",X"20",X"CD",X"48",X"16",
		X"D5",X"E5",X"3A",X"F8",X"4D",X"3C",X"32",X"F8",X"4D",X"FE",X"03",X"C2",X"2B",X"15",X"21",X"7E",
		X"1D",X"3A",X"F8",X"4D",X"CD",X"E3",X"15",X"7E",X"E1",X"D1",X"E5",X"CD",X"E8",X"15",X"21",X"F1",
		X"4D",X"01",X"03",X"00",X"ED",X"B0",X"3A",X"F8",X"4D",X"FE",X"00",X"28",X"25",X"21",X"82",X"1D",
		X"CD",X"E3",X"15",X"7E",X"D1",X"CD",X"52",X"16",X"21",X"F3",X"4D",X"CD",X"9C",X"11",X"21",X"B4",
		X"4D",X"11",X"F2",X"43",X"CD",X"ED",X"15",X"21",X"92",X"4D",X"CB",X"86",X"3E",X"01",X"CD",X"70",
		X"15",X"C9",X"D1",X"3E",X"80",X"CD",X"52",X"16",X"3E",X"20",X"CD",X"52",X"16",X"18",X"D9",X"3A",
		X"F7",X"4D",X"FE",X"00",X"CA",X"16",X"14",X"3D",X"32",X"F7",X"4D",X"FE",X"1A",X"28",X"14",X"3E",
		X"1B",X"2A",X"F9",X"4D",X"77",X"3E",X"20",X"CD",X"E3",X"15",X"22",X"F9",X"4D",X"3E",X"1A",X"77",
		X"C3",X"16",X"14",X"3D",X"32",X"F7",X"4D",X"3E",X"1B",X"2A",X"F9",X"4D",X"2B",X"77",X"23",X"77",
		X"23",X"77",X"2B",X"3E",X"40",X"18",X"E0",X"3A",X"F7",X"4D",X"FE",X"1B",X"CA",X"16",X"14",X"3C",
		X"32",X"F7",X"4D",X"FE",X"1A",X"28",X"14",X"3E",X"1B",X"2A",X"F9",X"4D",X"77",X"3E",X"20",X"CD",
		X"48",X"16",X"22",X"F9",X"4D",X"3E",X"1A",X"77",X"C3",X"16",X"14",X"3C",X"32",X"F7",X"4D",X"3E",
		X"1B",X"2A",X"F9",X"4D",X"77",X"3E",X"40",X"CD",X"48",X"16",X"22",X"F9",X"4D",X"3E",X"1A",X"2B",
		X"77",X"23",X"77",X"23",X"77",X"C3",X"16",X"14",X"3E",X"08",X"CD",X"CE",X"15",X"32",X"C0",X"50",
		X"06",X"14",X"CD",X"90",X"15",X"DA",X"4E",X"14",X"C3",X"FF",X"13",X"3A",X"F5",X"4D",X"21",X"92",
		X"4D",X"CB",X"66",X"28",X"03",X"3A",X"F6",X"4D",X"CB",X"67",X"32",X"C0",X"50",X"28",X"EC",X"18",
		X"DC",X"02",X"1B",X"18",X"1A",X"21",X"40",X"40",X"11",X"41",X"40",X"01",X"7F",X"03",X"77",X"ED",
		X"B0",X"32",X"C0",X"50",X"C9",X"21",X"40",X"44",X"11",X"41",X"44",X"01",X"7F",X"03",X"77",X"ED",
		X"B0",X"32",X"C0",X"50",X"C9",X"3E",X"02",X"CD",X"55",X"15",X"3E",X"40",X"CD",X"45",X"15",X"C9",
		X"47",X"AF",X"32",X"99",X"4D",X"32",X"9B",X"4D",X"3A",X"9B",X"4D",X"B8",X"C8",X"21",X"90",X"4D",
		X"CB",X"6E",X"C0",X"32",X"C0",X"50",X"18",X"F0",X"E5",X"21",X"20",X"00",X"19",X"EB",X"E1",X"C9",
		X"3A",X"92",X"4D",X"CB",X"47",X"28",X"0D",X"3A",X"9C",X"4D",X"47",X"3A",X"9B",X"4D",X"B8",X"30",
		X"19",X"37",X"3F",X"C9",X"78",X"32",X"9C",X"4D",X"3A",X"92",X"4D",X"CB",X"C7",X"32",X"92",X"4D",
		X"AF",X"32",X"9B",X"4D",X"32",X"99",X"4D",X"37",X"3F",X"C9",X"3A",X"92",X"4D",X"CB",X"87",X"32",
		X"92",X"4D",X"37",X"C9",X"21",X"90",X"4D",X"CB",X"FE",X"CB",X"7E",X"C8",X"18",X"FB",X"47",X"AF",
		X"32",X"9A",X"4D",X"3A",X"9A",X"4D",X"B8",X"C8",X"21",X"90",X"4D",X"CB",X"6E",X"C0",X"32",X"C0",
		X"50",X"18",X"F0",X"85",X"6F",X"D0",X"24",X"C9",X"83",X"5F",X"D0",X"14",X"C9",X"3E",X"03",X"F5",
		X"7E",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"3A",X"91",X"4D",X"CB",
		X"77",X"28",X"22",X"78",X"12",X"1B",X"7E",X"E6",X"0F",X"47",X"3A",X"91",X"4D",X"CB",X"77",X"32",
		X"91",X"4D",X"28",X"20",X"78",X"12",X"2B",X"1B",X"F1",X"3D",X"20",X"D3",X"3A",X"91",X"4D",X"CB",
		X"B7",X"32",X"91",X"4D",X"C9",X"78",X"FE",X"00",X"28",X"DB",X"3A",X"91",X"4D",X"CB",X"F7",X"32",
		X"91",X"4D",X"18",X"CF",X"78",X"FE",X"00",X"28",X"DD",X"3A",X"91",X"4D",X"CB",X"F7",X"32",X"91",
		X"4D",X"18",X"D1",X"81",X"4F",X"D0",X"04",X"C9",X"D5",X"16",X"00",X"5F",X"37",X"3F",X"ED",X"52",
		X"D1",X"C9",X"E5",X"EB",X"16",X"00",X"5F",X"37",X"3F",X"ED",X"52",X"EB",X"E1",X"C9",X"CD",X"5B",
		X"1A",X"DD",X"CB",X"00",X"D6",X"C9",X"32",X"F8",X"4C",X"D5",X"3A",X"F8",X"4C",X"4F",X"ED",X"A0",
		X"79",X"FE",X"00",X"20",X"F9",X"D1",X"CD",X"88",X"15",X"10",X"EE",X"C9",X"32",X"F8",X"4C",X"D5",
		X"3A",X"F8",X"4C",X"4F",X"ED",X"A0",X"2B",X"79",X"FE",X"00",X"20",X"F8",X"D1",X"CD",X"88",X"15",
		X"10",X"ED",X"C9",X"DD",X"7E",X"05",X"FD",X"96",X"05",X"B8",X"DA",X"E5",X"16",X"57",X"3E",X"FF",
		X"90",X"47",X"7A",X"B8",X"D2",X"E5",X"16",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"B9",X"DA",X"0F",
		X"17",X"57",X"3E",X"FF",X"91",X"4F",X"7A",X"B9",X"D2",X"0F",X"17",X"FD",X"7E",X"05",X"DD",X"BE",
		X"05",X"D2",X"24",X"17",X"FD",X"7E",X"04",X"DD",X"BE",X"04",X"D2",X"2C",X"17",X"3A",X"FF",X"4D",
		X"21",X"DD",X"16",X"CB",X"27",X"CD",X"E3",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"A9",X"17",X"82",
		X"17",X"34",X"17",X"5B",X"17",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"B9",X"38",X"18",X"57",X"3E",
		X"FF",X"91",X"4F",X"7A",X"B9",X"30",X"0F",X"DD",X"7E",X"04",X"FD",X"BE",X"04",X"38",X"0A",X"DD",
		X"36",X"00",X"18",X"3E",X"02",X"C9",X"3E",X"01",X"C9",X"DD",X"36",X"00",X"08",X"18",X"F4",X"DD",
		X"7E",X"05",X"FD",X"BE",X"05",X"38",X"07",X"DD",X"36",X"00",X"00",X"3E",X"03",X"C9",X"DD",X"36",
		X"00",X"10",X"18",X"F7",X"21",X"FF",X"4D",X"CB",X"C6",X"C3",X"C4",X"16",X"21",X"FF",X"4D",X"CB",
		X"CE",X"C3",X"CD",X"16",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"47",X"DD",X"7E",X"05",X"FD",X"96",
		X"05",X"B8",X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",X"02",X"C3",X"CD",X"17",X"DD",X"36",X"00",
		X"04",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"06",X"C3",X"CD",X"17",X"FD",X"7E",X"04",X"DD",X"96",
		X"04",X"47",X"FD",X"7E",X"05",X"DD",X"96",X"05",X"B8",X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",
		X"0E",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"0C",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"0A",X"C3",
		X"CD",X"17",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"47",X"FD",X"7E",X"05",X"DD",X"96",X"05",X"B8",
		X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",X"12",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"14",X"C3",
		X"CD",X"17",X"DD",X"36",X"00",X"16",X"C3",X"CD",X"17",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"47",
		X"DD",X"7E",X"05",X"FD",X"96",X"05",X"B8",X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",X"1E",X"C3",
		X"CD",X"17",X"DD",X"36",X"00",X"1C",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"1A",X"AF",X"32",X"FF",
		X"4D",X"C9",X"2A",X"FD",X"4D",X"E5",X"21",X"13",X"8C",X"7D",X"E1",X"BD",X"CC",X"0F",X"18",X"7E",
		X"FE",X"00",X"CA",X"F5",X"17",X"23",X"46",X"3A",X"75",X"4D",X"B8",X"CA",X"05",X"18",X"2B",X"22",
		X"FD",X"4D",X"C3",X"0E",X"18",X"23",X"46",X"3A",X"76",X"4D",X"B8",X"CA",X"05",X"18",X"2B",X"22",
		X"FD",X"4D",X"C3",X"0E",X"18",X"23",X"7E",X"32",X"F5",X"4D",X"23",X"22",X"FD",X"4D",X"C9",X"3E",
		X"FF",X"32",X"F5",X"4D",X"C9",X"3A",X"00",X"50",X"E6",X"0F",X"47",X"3A",X"40",X"50",X"E6",X"F0",
		X"B0",X"32",X"F5",X"4D",X"C9",X"3A",X"40",X"50",X"47",X"E6",X"0F",X"CB",X"78",X"28",X"02",X"CB",
		X"E7",X"32",X"F6",X"4D",X"C9",X"DD",X"21",X"02",X"4E",X"DD",X"CB",X"00",X"46",X"C4",X"5E",X"16",
		X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"51",X"50",X"CD",X"5E",X"19",
		X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"1D",X"4E",X"DD",X"CB",X"00",X"46",X"C4",X"5E",
		X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"51",X"50",X"CD",X"5E",
		X"19",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"38",X"4E",X"DD",X"CB",X"00",X"46",X"C4",
		X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"51",X"50",X"CD",
		X"5E",X"19",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"53",X"4E",X"DD",X"CB",X"00",X"46",
		X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"56",X"50",
		X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"6E",X"4E",X"DD",X"CB",X"00",
		X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"56",
		X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"89",X"4E",X"DD",X"CB",
		X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",
		X"56",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"A4",X"4E",X"DD",
		X"CB",X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",
		X"21",X"5B",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4F",X"50",X"DD",X"21",X"BF",X"4E",
		X"DD",X"CB",X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",
		X"FD",X"21",X"5B",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4F",X"50",X"DD",X"21",X"DA",
		X"4E",X"DD",X"CB",X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"C8",X"CD",X"87",X"19",
		X"FD",X"21",X"5B",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4F",X"50",X"C9",X"DD",X"7E",
		X"03",X"FD",X"77",X"00",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FD",X"77",X"01",X"DD",
		X"7E",X"04",X"FD",X"77",X"02",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FD",X"77",X"03",
		X"DD",X"7E",X"05",X"FD",X"77",X"04",X"C9",X"DD",X"CB",X"00",X"4E",X"C2",X"5B",X"1A",X"DD",X"6E",
		X"01",X"DD",X"66",X"02",X"7E",X"CB",X"27",X"11",X"A5",X"19",X"CD",X"E8",X"15",X"23",X"E5",X"1A",
		X"6F",X"13",X"1A",X"67",X"E9",X"BF",X"19",X"C3",X"19",X"D1",X"19",X"DA",X"19",X"F0",X"19",X"FD",
		X"19",X"17",X"1A",X"30",X"1A",X"52",X"1A",X"5A",X"1A",X"79",X"1A",X"85",X"1A",X"91",X"1A",X"E1",
		X"C3",X"94",X"19",X"E1",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"23",X"DD",X"77",X"04",X"C3",X"94",
		X"19",X"E1",X"7E",X"DD",X"77",X"05",X"23",X"C3",X"94",X"19",X"E1",X"7E",X"DD",X"46",X"03",X"80",
		X"DD",X"77",X"03",X"23",X"7E",X"23",X"DD",X"46",X"04",X"88",X"DD",X"77",X"04",X"C3",X"94",X"19",
		X"E1",X"7E",X"DD",X"46",X"05",X"80",X"DD",X"77",X"05",X"23",X"C3",X"94",X"19",X"E1",X"DD",X"7E",
		X"07",X"BE",X"30",X"0B",X"DD",X"34",X"07",X"2B",X"DD",X"75",X"01",X"DD",X"74",X"02",X"C9",X"DD",
		X"36",X"07",X"00",X"23",X"C3",X"94",X"19",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"D1",X"D5",X"2B",
		X"72",X"2B",X"73",X"2B",X"36",X"00",X"DD",X"75",X"08",X"DD",X"74",X"09",X"E1",X"C3",X"94",X"19",
		X"D1",X"1A",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"BE",X"28",X"09",X"34",X"23",X"5E",X"23",X"56",
		X"EB",X"C3",X"94",X"19",X"23",X"23",X"23",X"DD",X"75",X"08",X"DD",X"74",X"09",X"13",X"EB",X"C3",
		X"94",X"19",X"E1",X"5E",X"23",X"56",X"EB",X"C3",X"94",X"19",X"E1",X"DD",X"E5",X"DD",X"E5",X"E1",
		X"D1",X"13",X"36",X"00",X"01",X"18",X"00",X"ED",X"B0",X"1A",X"DD",X"77",X"01",X"13",X"1A",X"DD",
		X"77",X"02",X"DD",X"75",X"08",X"DD",X"74",X"09",X"C9",X"E1",X"DD",X"75",X"01",X"DD",X"74",X"02",
		X"DD",X"36",X"00",X"00",X"C9",X"E1",X"5E",X"23",X"56",X"EB",X"36",X"06",X"13",X"EB",X"C3",X"94",
		X"19",X"E1",X"7E",X"DD",X"77",X"06",X"23",X"C3",X"94",X"19",X"32",X"40",X"52",X"45",X"59",X"41",
		X"4C",X"50",X"40",X"45",X"52",X"4F",X"43",X"53",X"50",X"4F",X"54",X"40",X"31",X"40",X"52",X"45",
		X"59",X"41",X"4C",X"50",X"54",X"49",X"44",X"45",X"52",X"43",X"59",X"41",X"4C",X"50",X"45",X"45",
		X"52",X"46",X"40",X"4E",X"49",X"4F",X"43",X"40",X"54",X"52",X"45",X"53",X"4E",X"49",X"52",X"45",
		X"59",X"41",X"4C",X"50",X"40",X"45",X"4E",X"4F",X"40",X"54",X"43",X"45",X"4C",X"45",X"53",X"52",
		X"4F",X"53",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",X"4F",X"57",X"54",X"40",X"52",X"4F",X"40",
		X"45",X"4E",X"4F",X"40",X"54",X"43",X"45",X"4C",X"45",X"53",X"50",X"55",X"40",X"45",X"4E",X"4F",
		X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"50",X"55",X"40",X"4F",X"57",X"54",X"40",X"52",X"45",
		X"59",X"41",X"4C",X"50",X"52",X"45",X"56",X"4F",X"40",X"45",X"4D",X"41",X"47",X"59",X"52",X"44",
		X"52",X"41",X"5A",X"49",X"57",X"40",X"46",X"4F",X"40",X"4C",X"4C",X"41",X"48",X"45",X"48",X"54",
		X"40",X"4E",X"49",X"40",X"53",X"49",X"40",X"45",X"52",X"4F",X"43",X"53",X"40",X"52",X"55",X"4F",
		X"59",X"4E",X"45",X"54",X"40",X"50",X"4F",X"54",X"54",X"43",X"45",X"4C",X"45",X"53",X"40",X"4F",
		X"54",X"40",X"4B",X"43",X"49",X"54",X"53",X"59",X"4F",X"4A",X"40",X"45",X"53",X"55",X"4E",X"4F",
		X"54",X"54",X"55",X"42",X"40",X"45",X"52",X"49",X"46",X"40",X"44",X"4E",X"41",X"40",X"52",X"45",
		X"54",X"54",X"45",X"4C",X"54",X"4E",X"49",X"52",X"50",X"40",X"4F",X"54",X"45",X"4E",X"44",X"4D",
		X"41",X"4C",X"53",X"53",X"4E",X"4F",X"49",X"54",X"43",X"55",X"52",X"54",X"53",X"4E",X"49",X"40",
		X"59",X"41",X"4C",X"50",X"40",X"31",X"40",X"53",X"4E",X"49",X"4F",X"43",X"40",X"32",X"53",X"59",
		X"41",X"4C",X"50",X"40",X"32",X"40",X"40",X"4E",X"49",X"4F",X"43",X"40",X"31",X"40",X"59",X"41",
		X"4C",X"50",X"40",X"31",X"40",X"40",X"4E",X"49",X"4F",X"43",X"40",X"31",X"53",X"54",X"4E",X"49",
		X"4F",X"50",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"59",X"52",X"45",X"56",X"45",X"40",
		X"53",X"55",X"4E",X"4F",X"42",X"30",X"30",X"30",X"30",X"35",X"31",X"30",X"30",X"30",X"35",X"32",
		X"31",X"30",X"30",X"30",X"30",X"30",X"31",X"40",X"30",X"30",X"30",X"35",X"37",X"53",X"43",X"49",
		X"54",X"53",X"4F",X"4E",X"47",X"41",X"49",X"44",X"4E",X"4F",X"49",X"54",X"49",X"44",X"4E",X"4F",
		X"43",X"40",X"40",X"4E",X"4F",X"49",X"54",X"41",X"43",X"4F",X"4C",X"40",X"40",X"4D",X"4F",X"52",
		X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"44",X"37",X"40",X"40",X"40",
		X"40",X"40",X"40",X"31",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"46",
		X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"32",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"48",X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"33",X"44",X"4F",X"4F",X"47",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4A",X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"34",
		X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"48",X"34",X"40",X"40",X"40",
		X"40",X"40",X"40",X"31",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4C",
		X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"32",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"4A",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"33",X"44",X"4F",X"4F",X"47",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4D",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"34",
		X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4B",X"34",X"40",X"40",X"40",
		X"40",X"40",X"40",X"35",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4E",
		X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"36",X"44",X"41",X"42",X"40",X"4E",X"4F",X"49",X"54",
		X"49",X"44",X"4E",X"4F",X"43",X"40",X"40",X"4E",X"4F",X"49",X"54",X"41",X"43",X"4F",X"4C",X"40",
		X"40",X"4D",X"41",X"52",X"4E",X"45",X"4D",X"40",X"41",X"52",X"54",X"58",X"45",X"40",X"32",X"40",
		X"52",X"4F",X"46",X"06",X"03",X"1A",X"BE",X"38",X"08",X"20",X"0E",X"2B",X"1B",X"10",X"F6",X"18",
		X"06",X"CD",X"1E",X"1D",X"37",X"3F",X"C9",X"37",X"C9",X"CD",X"1E",X"1D",X"37",X"C9",X"78",X"FE",
		X"00",X"C8",X"2B",X"1B",X"3D",X"20",X"FB",X"C9",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",
		X"08",X"09",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",
		X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5A",X"59",X"58",X"57",
		X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"47",
		X"46",X"45",X"44",X"43",X"42",X"41",X"00",X"01",X"04",X"02",X"94",X"42",X"95",X"42",X"96",X"42",
		X"97",X"42",X"98",X"42",X"99",X"42",X"9A",X"42",X"9B",X"42",X"9C",X"42",X"9D",X"42",X"03",X"02",
		X"01",X"00",X"00",X"80",X"60",X"40",X"3A",X"FD",X"4E",X"A7",X"20",X"15",X"21",X"BF",X"4E",X"CB",
		X"56",X"28",X"0E",X"3A",X"2A",X"4F",X"3C",X"32",X"2A",X"4F",X"20",X"05",X"CB",X"CE",X"C3",X"11",
		X"31",X"3A",X"0B",X"4F",X"A7",X"C2",X"8C",X"30",X"21",X"09",X"4F",X"CB",X"7E",X"20",X"0E",X"35",
		X"20",X"0B",X"3A",X"53",X"4E",X"A7",X"28",X"05",X"CB",X"CF",X"32",X"53",X"4E",X"3A",X"77",X"4D",
		X"FE",X"78",X"DA",X"CA",X"1D",X"FE",X"90",X"DA",X"D7",X"1D",X"3A",X"5F",X"4D",X"FE",X"78",X"DA",
		X"0A",X"1E",X"FE",X"90",X"D2",X"0A",X"1E",X"3A",X"FE",X"4E",X"FE",X"01",X"C2",X"17",X"1E",X"3A",
		X"39",X"43",X"FE",X"E4",X"DA",X"F9",X"1D",X"3E",X"DD",X"32",X"39",X"43",X"32",X"F9",X"40",X"3C",
		X"32",X"19",X"43",X"32",X"D9",X"40",X"C3",X"17",X"1E",X"3E",X"E4",X"32",X"39",X"43",X"32",X"19",
		X"43",X"32",X"F9",X"40",X"32",X"D9",X"40",X"C3",X"17",X"1E",X"3A",X"39",X"43",X"FE",X"9A",X"CA",
		X"17",X"1E",X"3E",X"9A",X"C3",X"FB",X"1D",X"3A",X"80",X"4C",X"A7",X"CA",X"36",X"1E",X"DD",X"21",
		X"80",X"4C",X"21",X"A4",X"1E",X"3A",X"81",X"4C",X"A7",X"CA",X"58",X"1E",X"CD",X"6D",X"1E",X"DD",
		X"22",X"F4",X"4C",X"CD",X"16",X"0E",X"3A",X"90",X"4C",X"A7",X"CA",X"39",X"20",X"21",X"BC",X"1E",
		X"DD",X"21",X"90",X"4C",X"3A",X"91",X"4C",X"A7",X"CA",X"58",X"1E",X"CD",X"6D",X"1E",X"DD",X"22",
		X"F4",X"4C",X"CD",X"16",X"0E",X"C3",X"39",X"20",X"DD",X"36",X"01",X"10",X"DD",X"36",X"05",X"AE",
		X"DD",X"7E",X"09",X"CB",X"27",X"CD",X"E3",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"DD",X"7E",X"04",
		X"DD",X"96",X"08",X"C0",X"DD",X"7E",X"03",X"DD",X"96",X"07",X"CA",X"8A",X"1E",X"DA",X"85",X"1E",
		X"DD",X"36",X"00",X"04",X"C9",X"DD",X"36",X"00",X"05",X"C9",X"DD",X"36",X"00",X"00",X"DD",X"36",
		X"01",X"00",X"2A",X"8E",X"4D",X"CB",X"46",X"CA",X"9F",X"1E",X"DD",X"36",X"05",X"BE",X"C9",X"DD",
		X"36",X"05",X"BD",X"C9",X"D4",X"1E",X"E3",X"1E",X"F2",X"1E",X"01",X"1F",X"10",X"1F",X"1F",X"1F",
		X"2E",X"1F",X"3D",X"1F",X"4C",X"1F",X"5B",X"1F",X"6A",X"1F",X"79",X"1F",X"88",X"1F",X"97",X"1F",
		X"A6",X"1F",X"B5",X"1F",X"C4",X"1F",X"D3",X"1F",X"E2",X"1F",X"F1",X"1F",X"00",X"20",X"0F",X"20",
		X"1E",X"20",X"2D",X"20",X"DD",X"36",X"07",X"D0",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"01",
		X"C3",X"36",X"1E",X"DD",X"36",X"07",X"98",X"DD",X"36",X"08",X"E8",X"DD",X"36",X"09",X"02",X"C3",
		X"36",X"1E",X"DD",X"36",X"07",X"C8",X"DD",X"36",X"08",X"E8",X"DD",X"36",X"09",X"03",X"C3",X"36",
		X"1E",X"DD",X"36",X"07",X"D0",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"04",X"C3",X"36",X"1E",
		X"DD",X"36",X"07",X"A0",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"05",X"C3",X"36",X"1E",X"DD",
		X"36",X"07",X"A0",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"06",X"C3",X"36",X"1E",X"DD",X"36",
		X"07",X"D8",X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"07",X"C3",X"36",X"1E",X"DD",X"36",X"07",
		X"B8",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"08",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"A8",
		X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"09",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"C8",X"DD",
		X"36",X"08",X"F0",X"DD",X"36",X"09",X"0A",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"B0",X"DD",X"36",
		X"08",X"E8",X"DD",X"36",X"09",X"0B",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"B8",X"DD",X"36",X"08",
		X"E0",X"DD",X"36",X"09",X"0B",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"08",X"DD",X"36",X"08",X"F8",
		X"DD",X"36",X"09",X"01",X"C3",X"39",X"20",X"DD",X"36",X"07",X"40",X"DD",X"36",X"08",X"E8",X"DD",
		X"36",X"09",X"02",X"C3",X"39",X"20",X"DD",X"36",X"07",X"10",X"DD",X"36",X"08",X"E8",X"DD",X"36",
		X"09",X"03",X"C3",X"39",X"20",X"DD",X"36",X"07",X"08",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",
		X"04",X"C3",X"39",X"20",X"DD",X"36",X"07",X"38",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"05",
		X"C3",X"39",X"20",X"DD",X"36",X"07",X"38",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"06",X"C3",
		X"39",X"20",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"07",X"C3",X"39",
		X"20",X"DD",X"36",X"07",X"20",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"08",X"C3",X"39",X"20",
		X"DD",X"36",X"07",X"30",X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"09",X"C3",X"39",X"20",X"DD",
		X"36",X"07",X"10",X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"0A",X"C3",X"39",X"20",X"DD",X"36",
		X"07",X"28",X"DD",X"36",X"08",X"E8",X"DD",X"36",X"09",X"0B",X"C3",X"39",X"20",X"DD",X"36",X"07",
		X"20",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"0B",X"3A",X"91",X"4D",X"CB",X"6F",X"28",X"16",
		X"DD",X"21",X"71",X"4D",X"AF",X"32",X"22",X"4F",X"3A",X"F5",X"4D",X"32",X"23",X"4F",X"CD",X"D2",
		X"2F",X"3A",X"0B",X"4F",X"A7",X"C0",X"3A",X"91",X"4D",X"CB",X"4F",X"28",X"17",X"DD",X"21",X"59",
		X"4D",X"3E",X"01",X"32",X"22",X"4F",X"3A",X"F6",X"4D",X"32",X"23",X"4F",X"CD",X"D2",X"2F",X"3A",
		X"0B",X"4F",X"A7",X"C0",X"21",X"FF",X"4E",X"34",X"20",X"43",X"21",X"00",X"4F",X"34",X"46",X"3A",
		X"08",X"4F",X"B8",X"20",X"38",X"21",X"FF",X"4E",X"35",X"35",X"23",X"35",X"3A",X"24",X"4D",X"FE",
		X"50",X"38",X"2A",X"CB",X"7F",X"20",X"22",X"DD",X"21",X"11",X"4D",X"CD",X"71",X"26",X"3A",X"15",
		X"4D",X"A7",X"28",X"19",X"DD",X"36",X"13",X"0A",X"3A",X"17",X"4D",X"C6",X"18",X"32",X"17",X"4D",
		X"21",X"BF",X"4E",X"CB",X"C6",X"DD",X"21",X"59",X"4D",X"AF",X"32",X"00",X"4F",X"3A",X"FF",X"4E",
		X"CB",X"47",X"28",X"04",X"DD",X"21",X"71",X"4D",X"DD",X"7E",X"0B",X"32",X"FD",X"4C",X"DD",X"7E",
		X"0C",X"32",X"FE",X"4C",X"DD",X"7E",X"0D",X"32",X"FF",X"4C",X"21",X"FE",X"4E",X"35",X"20",X"06",
		X"36",X"06",X"21",X"01",X"4F",X"34",X"3A",X"25",X"4F",X"A7",X"C2",X"E2",X"2C",X"21",X"FA",X"4E",
		X"35",X"C2",X"10",X"21",X"DD",X"21",X"41",X"4D",X"2B",X"7E",X"3C",X"E6",X"F3",X"77",X"3A",X"54",
		X"4D",X"FE",X"20",X"D2",X"EA",X"21",X"CD",X"8E",X"2A",X"DD",X"36",X"0F",X"01",X"C3",X"D2",X"22",
		X"7E",X"FE",X"02",X"CA",X"9F",X"22",X"DA",X"D4",X"21",X"FE",X"BF",X"CA",X"7B",X"21",X"FE",X"BC",
		X"CA",X"9F",X"22",X"FE",X"04",X"30",X"32",X"3A",X"24",X"4D",X"FE",X"20",X"D2",X"59",X"21",X"DD",
		X"21",X"11",X"4D",X"CD",X"8E",X"2A",X"DD",X"36",X"0F",X"01",X"DD",X"36",X"01",X"18",X"DD",X"36",
		X"08",X"50",X"3A",X"15",X"4D",X"FE",X"01",X"C2",X"D2",X"22",X"DD",X"36",X"00",X"18",X"DD",X"36",
		X"04",X"FF",X"DD",X"36",X"06",X"24",X"C3",X"D2",X"22",X"3A",X"2D",X"4D",X"A7",X"C2",X"6A",X"21",
		X"DD",X"21",X"29",X"4D",X"CD",X"71",X"26",X"C3",X"EA",X"21",X"3A",X"45",X"4D",X"A7",X"C2",X"EA",
		X"21",X"DD",X"21",X"41",X"4D",X"CD",X"71",X"26",X"C3",X"EA",X"21",X"3A",X"91",X"4D",X"CB",X"6F",
		X"28",X"3B",X"3A",X"79",X"4D",X"E6",X"30",X"C2",X"BD",X"21",X"DD",X"21",X"71",X"4D",X"FD",X"21",
		X"29",X"4D",X"01",X"30",X"50",X"CD",X"66",X"04",X"DA",X"B5",X"21",X"FD",X"21",X"41",X"4D",X"01",
		X"30",X"50",X"CD",X"66",X"04",X"DA",X"B5",X"21",X"DD",X"36",X"06",X"74",X"DD",X"CB",X"08",X"E6",
		X"21",X"A4",X"4E",X"CB",X"C6",X"3E",X"C0",X"32",X"FA",X"4E",X"C3",X"D2",X"22",X"3A",X"91",X"4D",
		X"CB",X"4F",X"CA",X"EA",X"21",X"3A",X"61",X"4D",X"E6",X"30",X"C2",X"EA",X"21",X"DD",X"21",X"59",
		X"4D",X"C3",X"8E",X"21",X"DD",X"21",X"29",X"4D",X"3A",X"3C",X"4D",X"FE",X"20",X"D2",X"EA",X"21",
		X"CD",X"8E",X"2A",X"DD",X"36",X"0F",X"01",X"C3",X"D2",X"22",X"DD",X"21",X"29",X"4D",X"3A",X"3C",
		X"4D",X"FE",X"20",X"D2",X"FD",X"21",X"21",X"38",X"4D",X"35",X"CA",X"F8",X"23",X"DD",X"21",X"41",
		X"4D",X"3A",X"54",X"4D",X"FE",X"20",X"D2",X"10",X"22",X"21",X"50",X"4D",X"35",X"CA",X"F8",X"23",
		X"DD",X"21",X"11",X"4D",X"3A",X"24",X"4D",X"FE",X"20",X"D2",X"23",X"22",X"21",X"20",X"4D",X"35",
		X"CA",X"F8",X"23",X"DD",X"21",X"29",X"4D",X"3A",X"3C",X"4D",X"CB",X"7F",X"C2",X"D2",X"22",X"FE",
		X"40",X"D2",X"3B",X"22",X"21",X"31",X"4D",X"35",X"CA",X"BB",X"24",X"DD",X"21",X"41",X"4D",X"3A",
		X"54",X"4D",X"CB",X"7F",X"C2",X"D2",X"22",X"FE",X"40",X"D2",X"53",X"22",X"21",X"49",X"4D",X"35",
		X"CA",X"BB",X"24",X"DD",X"21",X"11",X"4D",X"3A",X"24",X"4D",X"CB",X"7F",X"C2",X"D2",X"22",X"FE",
		X"40",X"D2",X"D2",X"22",X"21",X"19",X"4D",X"35",X"CA",X"BB",X"24",X"C3",X"D2",X"22",X"91",X"4C",
		X"49",X"5A",X"41",X"52",X"44",X"20",X"57",X"49",X"5A",X"41",X"52",X"44",X"2C",X"43",X"4F",X"50",
		X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"54",X"45",X"43",X"48",X"53",
		X"54",X"41",X"52",X"20",X"49",X"4E",X"43",X"2E",X"DD",X"21",X"29",X"4D",X"C3",X"B6",X"22",X"3A",
		X"3C",X"4D",X"E6",X"70",X"FE",X"50",X"28",X"F0",X"3A",X"54",X"4D",X"E6",X"70",X"FE",X"50",X"C2",
		X"EA",X"21",X"DD",X"21",X"41",X"4D",X"DD",X"36",X"13",X"0A",X"DD",X"36",X"0F",X"08",X"DD",X"36",
		X"01",X"10",X"DD",X"7E",X"04",X"FE",X"01",X"20",X"04",X"DD",X"36",X"04",X"FF",X"3E",X"18",X"32",
		X"FA",X"4E",X"3A",X"FD",X"4E",X"FE",X"32",X"D4",X"DD",X"2C",X"FE",X"01",X"CA",X"BB",X"23",X"D2",
		X"A3",X"23",X"3A",X"77",X"4D",X"FE",X"90",X"30",X"05",X"FE",X"78",X"D2",X"A3",X"23",X"3A",X"5F",
		X"4D",X"FE",X"90",X"30",X"05",X"FE",X"78",X"D2",X"A3",X"23",X"3E",X"80",X"32",X"19",X"4D",X"32",
		X"31",X"4D",X"32",X"49",X"4D",X"3A",X"3C",X"4D",X"CB",X"7F",X"C2",X"A3",X"23",X"3A",X"54",X"4D",
		X"CB",X"7F",X"C2",X"A3",X"23",X"3A",X"24",X"4D",X"CB",X"7F",X"C2",X"A3",X"23",X"3A",X"3C",X"4D",
		X"FE",X"40",X"30",X"09",X"AF",X"32",X"2A",X"4D",X"3E",X"5A",X"32",X"3C",X"4D",X"3A",X"54",X"4D",
		X"FE",X"40",X"30",X"09",X"AF",X"32",X"42",X"4D",X"3E",X"5A",X"32",X"54",X"4D",X"3A",X"24",X"4D",
		X"FE",X"40",X"30",X"09",X"AF",X"32",X"12",X"4D",X"3E",X"5A",X"32",X"24",X"4D",X"3A",X"76",X"4D",
		X"FE",X"C9",X"30",X"4F",X"3A",X"5E",X"4D",X"FE",X"C9",X"30",X"48",X"3A",X"79",X"4D",X"CB",X"7F",
		X"28",X"41",X"E6",X"CF",X"32",X"79",X"4D",X"AF",X"32",X"FA",X"4E",X"3A",X"61",X"4D",X"CB",X"7F",
		X"28",X"31",X"E6",X"CF",X"32",X"61",X"4D",X"AF",X"32",X"5A",X"4D",X"32",X"72",X"4D",X"3A",X"53",
		X"4E",X"CB",X"4F",X"20",X"03",X"A7",X"20",X"1B",X"3A",X"81",X"4C",X"A7",X"20",X"15",X"3A",X"91",
		X"4C",X"A7",X"20",X"0F",X"3A",X"7E",X"4D",X"FE",X"90",X"20",X"08",X"3A",X"66",X"4D",X"FE",X"90",
		X"CA",X"61",X"30",X"DD",X"21",X"29",X"4D",X"CD",X"79",X"25",X"DD",X"21",X"41",X"4D",X"CD",X"79",
		X"25",X"DD",X"21",X"11",X"4D",X"CD",X"79",X"25",X"C3",X"4A",X"2C",X"3A",X"3C",X"4D",X"47",X"E6",
		X"0F",X"FE",X"0A",X"30",X"13",X"78",X"E6",X"70",X"FE",X"30",X"28",X"0C",X"78",X"E6",X"F0",X"F6",
		X"0A",X"32",X"3C",X"4D",X"AF",X"32",X"F8",X"4E",X"3A",X"54",X"4D",X"47",X"E6",X"0F",X"FE",X"0A",
		X"30",X"C1",X"78",X"E6",X"70",X"FE",X"30",X"28",X"BA",X"78",X"E6",X"F0",X"F6",X"0A",X"32",X"54",
		X"4D",X"AF",X"32",X"F8",X"4E",X"C3",X"A3",X"23",X"DD",X"7E",X"10",X"DD",X"77",X"0F",X"DD",X"7E",
		X"13",X"E6",X"0F",X"FE",X"0E",X"CA",X"0E",X"24",X"D2",X"58",X"24",X"C3",X"23",X"22",X"FD",X"21",
		X"71",X"4D",X"FD",X"CB",X"08",X"66",X"CA",X"58",X"24",X"01",X"00",X"00",X"CD",X"93",X"16",X"3A",
		X"FC",X"4D",X"FE",X"00",X"30",X"15",X"DD",X"7E",X"07",X"FE",X"08",X"28",X"0E",X"DD",X"7E",X"00",
		X"C6",X"10",X"FE",X"20",X"38",X"02",X"D6",X"20",X"DD",X"77",X"00",X"DD",X"7E",X"00",X"FE",X"10",
		X"CA",X"D2",X"22",X"D2",X"51",X"24",X"A7",X"CA",X"D2",X"22",X"DD",X"CB",X"06",X"CE",X"C3",X"D2",
		X"22",X"DD",X"CB",X"06",X"8E",X"C3",X"D2",X"22",X"FD",X"21",X"59",X"4D",X"FD",X"CB",X"08",X"66",
		X"CA",X"9B",X"24",X"01",X"00",X"00",X"CD",X"93",X"16",X"3A",X"FC",X"4D",X"FE",X"00",X"30",X"15",
		X"DD",X"7E",X"07",X"FE",X"08",X"28",X"0E",X"DD",X"7E",X"00",X"C6",X"10",X"FE",X"20",X"38",X"02",
		X"D6",X"20",X"DD",X"77",X"00",X"DD",X"7E",X"00",X"FE",X"10",X"CA",X"D2",X"22",X"D2",X"A6",X"24",
		X"A7",X"CA",X"D2",X"22",X"DD",X"CB",X"06",X"CE",X"C3",X"D2",X"22",X"3A",X"79",X"4D",X"CB",X"67",
		X"C2",X"0E",X"24",X"C3",X"D2",X"22",X"DD",X"CB",X"06",X"8E",X"C3",X"D2",X"22",X"DD",X"CB",X"07",
		X"5E",X"CA",X"23",X"22",X"DD",X"36",X"08",X"01",X"C3",X"D2",X"22",X"DD",X"36",X"08",X"03",X"DD",
		X"7E",X"05",X"E6",X"07",X"C2",X"AD",X"24",X"DD",X"7E",X"04",X"47",X"3E",X"F0",X"90",X"32",X"F3",
		X"4C",X"DD",X"7E",X"05",X"D6",X"10",X"32",X"F2",X"4C",X"CD",X"D0",X"0D",X"21",X"20",X"00",X"19",
		X"DD",X"7E",X"06",X"CB",X"4F",X"3A",X"A1",X"4C",X"C2",X"F6",X"24",X"FE",X"04",X"D2",X"AD",X"24",
		X"11",X"20",X"00",X"C3",X"FE",X"24",X"FE",X"05",X"DA",X"AD",X"24",X"11",X"E0",X"FF",X"DD",X"7E",
		X"0D",X"A7",X"C2",X"0E",X"25",X"3A",X"F7",X"4E",X"DD",X"77",X"08",X"C3",X"D2",X"22",X"47",X"4F",
		X"DD",X"75",X"09",X"DD",X"74",X"0A",X"19",X"7E",X"FE",X"9A",X"C2",X"6B",X"25",X"10",X"F7",X"DD",
		X"71",X"11",X"3A",X"F7",X"4E",X"DD",X"77",X"08",X"DD",X"36",X"01",X"00",X"DD",X"36",X"0B",X"CD",
		X"DD",X"CB",X"13",X"FE",X"DD",X"7E",X"06",X"FE",X"18",X"DA",X"4B",X"25",X"FE",X"30",X"DA",X"59",
		X"25",X"E6",X"03",X"C6",X"58",X"DD",X"77",X"06",X"C3",X"D2",X"22",X"E6",X"03",X"C6",X"14",X"DD",
		X"77",X"06",X"DD",X"CB",X"13",X"E6",X"C3",X"D2",X"22",X"E6",X"03",X"C6",X"2C",X"DD",X"77",X"06",
		X"DD",X"36",X"08",X"55",X"DD",X"CB",X"13",X"E6",X"C3",X"D2",X"22",X"FE",X"CD",X"DA",X"D2",X"22",
		X"79",X"90",X"CA",X"D2",X"22",X"4F",X"C3",X"1F",X"25",X"DD",X"7E",X"13",X"E6",X"70",X"FE",X"10",
		X"CA",X"13",X"27",X"DA",X"EA",X"27",X"FE",X"30",X"CA",X"94",X"25",X"DA",X"D6",X"26",X"FE",X"40",
		X"CA",X"33",X"26",X"C9",X"3A",X"FE",X"4E",X"FE",X"01",X"C2",X"13",X"2A",X"DD",X"36",X"01",X"10",
		X"DD",X"7E",X"0D",X"FE",X"07",X"30",X"06",X"DD",X"34",X"0D",X"DD",X"34",X"0D",X"3E",X"F0",X"DD",
		X"86",X"10",X"FE",X"0F",X"38",X"03",X"DD",X"77",X"10",X"3E",X"02",X"32",X"FA",X"4E",X"DD",X"7E",
		X"06",X"D6",X"14",X"DD",X"77",X"06",X"DD",X"7E",X"13",X"E6",X"0F",X"FE",X"04",X"DD",X"36",X"13",
		X"0A",X"CA",X"07",X"26",X"D2",X"10",X"26",X"FE",X"02",X"CA",X"F5",X"25",X"D2",X"FE",X"25",X"A7",
		X"C2",X"EC",X"25",X"21",X"00",X"4C",X"CD",X"96",X"3A",X"C3",X"13",X"2A",X"21",X"10",X"4C",X"CD",
		X"96",X"3A",X"C3",X"13",X"2A",X"21",X"20",X"4C",X"CD",X"96",X"3A",X"C3",X"13",X"2A",X"21",X"30",
		X"4C",X"CD",X"96",X"3A",X"C3",X"13",X"2A",X"21",X"40",X"4C",X"CD",X"96",X"3A",X"C3",X"13",X"2A",
		X"FE",X"06",X"CA",X"21",X"26",X"D2",X"2A",X"26",X"21",X"50",X"4C",X"CD",X"96",X"3A",X"C3",X"13",
		X"2A",X"21",X"60",X"4C",X"CD",X"96",X"3A",X"C3",X"13",X"2A",X"21",X"70",X"4C",X"CD",X"96",X"3A",
		X"C3",X"13",X"2A",X"DD",X"CB",X"13",X"7E",X"C2",X"61",X"26",X"CD",X"41",X"26",X"D0",X"C3",X"71",
		X"26",X"DD",X"7E",X"05",X"FE",X"05",X"D8",X"3A",X"FE",X"4E",X"FE",X"01",X"C0",X"DD",X"7E",X"06",
		X"47",X"E6",X"FC",X"4F",X"04",X"78",X"E6",X"03",X"81",X"DD",X"77",X"06",X"DD",X"36",X"01",X"20",
		X"C9",X"DD",X"7E",X"0B",X"FE",X"9A",X"CA",X"1B",X"27",X"3E",X"D0",X"DD",X"77",X"0B",X"C3",X"7A",
		X"27",X"DD",X"36",X"01",X"00",X"2A",X"8E",X"4D",X"7E",X"E6",X"07",X"FE",X"02",X"CA",X"BE",X"26",
		X"DA",X"CA",X"26",X"FE",X"03",X"CA",X"B2",X"26",X"11",X"91",X"40",X"21",X"01",X"88",X"01",X"18",
		X"0C",X"1A",X"FE",X"D3",X"C0",X"DD",X"71",X"00",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"70",
		X"06",X"DD",X"36",X"0F",X"01",X"DD",X"7E",X"13",X"E6",X"70",X"FE",X"60",X"C8",X"DD",X"36",X"13",
		X"5A",X"C9",X"11",X"51",X"43",X"21",X"0F",X"88",X"01",X"08",X"0E",X"C3",X"91",X"26",X"11",X"87",
		X"40",X"21",X"01",X"38",X"01",X"18",X"0C",X"C3",X"91",X"26",X"11",X"47",X"43",X"21",X"0F",X"38",
		X"01",X"08",X"0E",X"C3",X"91",X"26",X"DD",X"7E",X"05",X"FE",X"11",X"D2",X"0C",X"27",X"DD",X"7E",
		X"06",X"E6",X"03",X"C6",X"20",X"DD",X"77",X"06",X"DD",X"36",X"00",X"10",X"DD",X"36",X"01",X"15",
		X"DD",X"36",X"07",X"14",X"DD",X"36",X"0D",X"07",X"3E",X"02",X"32",X"FA",X"4E",X"DD",X"36",X"10",
		X"0F",X"DD",X"36",X"12",X"00",X"DD",X"36",X"13",X"0A",X"C3",X"13",X"2A",X"DD",X"CB",X"13",X"7E",
		X"CA",X"F3",X"27",X"DD",X"7E",X"0B",X"FE",X"9A",X"C2",X"7A",X"27",X"DD",X"35",X"11",X"FA",X"43",
		X"27",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"DD",X"CB",X"06",X"4E",X"CA",X"3D",X"27",X"01",X"20",
		X"00",X"36",X"9A",X"09",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"C3",X"13",X"2A",X"01",X"E0",X"FF",
		X"C3",X"31",X"27",X"DD",X"7E",X"06",X"D6",X"0C",X"DD",X"77",X"06",X"DD",X"36",X"0F",X"01",X"DD",
		X"36",X"01",X"10",X"FE",X"30",X"DD",X"CB",X"13",X"BE",X"D2",X"13",X"2A",X"DD",X"CB",X"13",X"A6",
		X"FE",X"18",X"DA",X"88",X"28",X"DD",X"CB",X"07",X"5E",X"C2",X"73",X"27",X"DD",X"36",X"01",X"15",
		X"C3",X"13",X"2A",X"DD",X"36",X"01",X"18",X"C3",X"13",X"2A",X"DD",X"7E",X"11",X"47",X"DD",X"7E",
		X"0C",X"90",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"CA",X"B4",X"27",X"DD",X"34",X"0C",X"DD",X"CB",
		X"06",X"4E",X"DD",X"7E",X"0B",X"CA",X"A6",X"27",X"01",X"E0",X"FF",X"09",X"77",X"DD",X"75",X"09",
		X"DD",X"74",X"0A",X"C3",X"13",X"2A",X"01",X"20",X"00",X"09",X"77",X"DD",X"75",X"09",X"DD",X"74",
		X"0A",X"C3",X"13",X"2A",X"DD",X"7E",X"0B",X"FE",X"D0",X"CA",X"DF",X"27",X"DD",X"34",X"0B",X"DD",
		X"CB",X"06",X"4E",X"CA",X"D9",X"27",X"11",X"20",X"00",X"19",X"10",X"FD",X"DD",X"75",X"09",X"DD",
		X"74",X"0A",X"DD",X"36",X"0C",X"00",X"C3",X"13",X"2A",X"11",X"E0",X"FF",X"C3",X"C9",X"27",X"DD",
		X"36",X"0B",X"9A",X"DD",X"36",X"0C",X"00",X"C3",X"13",X"2A",X"CD",X"B1",X"3A",X"D2",X"F3",X"27",
		X"DD",X"34",X"12",X"3A",X"FE",X"4E",X"FE",X"06",X"28",X"05",X"FE",X"03",X"C2",X"88",X"28",X"DD",
		X"7E",X"06",X"47",X"E6",X"FC",X"FE",X"58",X"DA",X"21",X"28",X"FE",X"5C",X"C2",X"18",X"28",X"78",
		X"C6",X"FC",X"DD",X"77",X"06",X"C3",X"13",X"2A",X"78",X"C6",X"04",X"DD",X"77",X"06",X"C3",X"13",
		X"2A",X"DD",X"CB",X"12",X"46",X"CA",X"5C",X"28",X"DD",X"35",X"05",X"78",X"E6",X"FC",X"FE",X"30",
		X"DA",X"3D",X"28",X"C2",X"0F",X"28",X"DD",X"CB",X"12",X"86",X"C3",X"18",X"28",X"FE",X"18",X"CA",
		X"4F",X"28",X"A7",X"CA",X"4F",X"28",X"78",X"C6",X"FC",X"DD",X"77",X"06",X"C3",X"88",X"28",X"DD",
		X"CB",X"12",X"86",X"78",X"C6",X"04",X"DD",X"77",X"06",X"C3",X"88",X"28",X"DD",X"34",X"05",X"78",
		X"E6",X"FC",X"FE",X"10",X"DA",X"53",X"28",X"CA",X"7E",X"28",X"FE",X"28",X"DA",X"53",X"28",X"CA",
		X"7E",X"28",X"FE",X"54",X"DA",X"18",X"28",X"DD",X"CB",X"12",X"C6",X"C3",X"0F",X"28",X"DD",X"CB",
		X"12",X"C6",X"78",X"C6",X"FC",X"DD",X"77",X"06",X"DD",X"7E",X"13",X"FE",X"20",X"D2",X"13",X"2A",
		X"E6",X"0F",X"FE",X"0A",X"D2",X"13",X"2A",X"4F",X"FE",X"03",X"CA",X"2A",X"29",X"D2",X"AE",X"28",
		X"FE",X"01",X"CA",X"30",X"29",X"D2",X"24",X"29",X"21",X"03",X"4C",X"C3",X"15",X"29",X"FE",X"06",
		X"CA",X"36",X"29",X"D2",X"3C",X"29",X"FE",X"04",X"CA",X"12",X"29",X"21",X"53",X"4C",X"C3",X"15",
		X"29",X"3E",X"F0",X"DD",X"86",X"05",X"47",X"DD",X"CB",X"06",X"4E",X"C2",X"42",X"29",X"AF",X"DD",
		X"96",X"04",X"BB",X"CA",X"07",X"29",X"DA",X"F0",X"28",X"78",X"C6",X"05",X"92",X"DA",X"52",X"29",
		X"FE",X"0A",X"DA",X"47",X"29",X"DD",X"36",X"00",X"04",X"DD",X"CB",X"06",X"CE",X"C3",X"13",X"2A",
		X"78",X"C6",X"05",X"92",X"DA",X"68",X"29",X"FE",X"0A",X"DA",X"5D",X"29",X"DD",X"36",X"00",X"1C",
		X"DD",X"CB",X"06",X"8E",X"C3",X"13",X"2A",X"78",X"BA",X"DA",X"73",X"29",X"C2",X"7A",X"29",X"C3",
		X"81",X"29",X"21",X"43",X"4C",X"5E",X"23",X"56",X"23",X"7E",X"FE",X"AD",X"DA",X"C1",X"28",X"3E",
		X"F8",X"C3",X"C3",X"28",X"21",X"23",X"4C",X"C3",X"15",X"29",X"21",X"33",X"4C",X"C3",X"15",X"29",
		X"21",X"13",X"4C",X"C3",X"15",X"29",X"21",X"63",X"4C",X"C3",X"15",X"29",X"21",X"73",X"4C",X"C3",
		X"15",X"29",X"3E",X"E8",X"C3",X"CF",X"28",X"DD",X"36",X"00",X"08",X"DD",X"CB",X"06",X"CE",X"C3",
		X"13",X"2A",X"DD",X"36",X"00",X"0C",X"DD",X"CB",X"06",X"CE",X"C3",X"13",X"2A",X"DD",X"36",X"00",
		X"18",X"DD",X"CB",X"06",X"8E",X"C3",X"13",X"2A",X"DD",X"36",X"00",X"14",X"DD",X"CB",X"06",X"8E",
		X"C3",X"13",X"2A",X"DD",X"36",X"00",X"10",X"C3",X"13",X"2A",X"DD",X"36",X"00",X"00",X"C3",X"13",
		X"2A",X"7E",X"FE",X"AD",X"DA",X"FD",X"29",X"21",X"F8",X"4E",X"79",X"FE",X"03",X"CA",X"A3",X"29",
		X"D2",X"BB",X"29",X"FE",X"01",X"CA",X"AB",X"29",X"D2",X"B3",X"29",X"CB",X"86",X"21",X"00",X"4C",
		X"C3",X"E5",X"29",X"CB",X"9E",X"21",X"30",X"4C",X"C3",X"E5",X"29",X"CB",X"8E",X"21",X"10",X"4C",
		X"C3",X"E5",X"29",X"CB",X"96",X"21",X"20",X"4C",X"C3",X"E5",X"29",X"FE",X"06",X"CA",X"D0",X"29",
		X"D2",X"D8",X"29",X"FE",X"04",X"CA",X"E0",X"29",X"CB",X"AE",X"21",X"50",X"4C",X"C3",X"E5",X"29",
		X"CB",X"B6",X"21",X"60",X"4C",X"C3",X"E5",X"29",X"CB",X"BE",X"21",X"70",X"4C",X"C3",X"E5",X"29",
		X"CB",X"A6",X"21",X"40",X"4C",X"CD",X"96",X"3A",X"DD",X"36",X"00",X"00",X"DD",X"7E",X"06",X"E6",
		X"03",X"C6",X"38",X"DD",X"77",X"06",X"DD",X"36",X"13",X"2A",X"C3",X"13",X"2A",X"DD",X"7E",X"06",
		X"E6",X"03",X"C6",X"14",X"DD",X"77",X"06",X"DD",X"CB",X"13",X"E6",X"DD",X"CB",X"13",X"EE",X"DD",
		X"36",X"01",X"00",X"DD",X"7E",X"13",X"E6",X"70",X"FE",X"40",X"D0",X"3A",X"79",X"4D",X"E6",X"30",
		X"FE",X"10",X"20",X"54",X"FD",X"21",X"71",X"4D",X"01",X"08",X"08",X"CD",X"66",X"04",X"30",X"48",
		X"FD",X"7E",X"08",X"E6",X"C0",X"F6",X"26",X"FD",X"77",X"08",X"FD",X"36",X"00",X"10",X"CD",X"F4",
		X"2A",X"DD",X"7E",X"13",X"E6",X"80",X"F6",X"4A",X"DD",X"77",X"13",X"DD",X"36",X"01",X"20",X"DD",
		X"36",X"00",X"10",X"FD",X"7E",X"04",X"FD",X"77",X"0B",X"FD",X"7E",X"05",X"FD",X"77",X"0C",X"FD",
		X"36",X"0D",X"98",X"FD",X"36",X"17",X"90",X"21",X"53",X"4E",X"CB",X"C6",X"DD",X"7E",X"07",X"FE",
		X"08",X"C0",X"21",X"A4",X"4E",X"CB",X"C6",X"C9",X"3A",X"61",X"4D",X"E6",X"30",X"FE",X"10",X"C0",
		X"FD",X"21",X"59",X"4D",X"01",X"08",X"08",X"CD",X"66",X"04",X"D0",X"C3",X"30",X"2A",X"3A",X"79",
		X"4D",X"CB",X"67",X"C2",X"B3",X"2A",X"3A",X"61",X"4D",X"CB",X"67",X"C2",X"B3",X"2A",X"3E",X"C0",
		X"32",X"FA",X"4E",X"DD",X"CB",X"06",X"4E",X"20",X"05",X"DD",X"36",X"00",X"1C",X"C9",X"DD",X"36",
		X"00",X"04",X"C9",X"DD",X"7E",X"06",X"FE",X"18",X"D2",X"21",X"2C",X"3A",X"F9",X"4E",X"CB",X"47",
		X"CA",X"21",X"2C",X"3A",X"F8",X"4E",X"FE",X"10",X"DA",X"DD",X"2A",X"CB",X"7F",X"C2",X"60",X"2B",
		X"CB",X"77",X"C2",X"73",X"2B",X"CB",X"6F",X"C2",X"86",X"2B",X"C3",X"99",X"2B",X"CB",X"5F",X"C2",
		X"AC",X"2B",X"CB",X"57",X"C2",X"BF",X"2B",X"CB",X"4F",X"C2",X"D2",X"2B",X"CB",X"47",X"C2",X"E5",
		X"2B",X"C3",X"21",X"2C",X"DD",X"7E",X"13",X"E6",X"0F",X"FE",X"0A",X"D0",X"FE",X"03",X"CA",X"45",
		X"2B",X"D2",X"15",X"2B",X"FE",X"01",X"CA",X"57",X"2B",X"D2",X"4E",X"2B",X"3A",X"F8",X"4E",X"CB",
		X"C7",X"32",X"F8",X"4E",X"C9",X"FE",X"06",X"CA",X"33",X"2B",X"D2",X"2A",X"2B",X"FE",X"04",X"28",
		X"1B",X"3A",X"F8",X"4E",X"CB",X"EF",X"32",X"F8",X"4E",X"C9",X"3A",X"F8",X"4E",X"CB",X"FF",X"32",
		X"F8",X"4E",X"C9",X"3A",X"F8",X"4E",X"CB",X"F7",X"32",X"F8",X"4E",X"C9",X"3A",X"F8",X"4E",X"CB",
		X"E7",X"32",X"F8",X"4E",X"C9",X"3A",X"F8",X"4E",X"CB",X"DF",X"32",X"F8",X"4E",X"C9",X"3A",X"F8",
		X"4E",X"CB",X"D7",X"32",X"F8",X"4E",X"C9",X"3A",X"F8",X"4E",X"CB",X"CF",X"32",X"F8",X"4E",X"C9",
		X"3A",X"73",X"4C",X"57",X"1E",X"07",X"CD",X"F8",X"2B",X"D0",X"3A",X"F8",X"4E",X"CB",X"BF",X"32",
		X"F8",X"4E",X"C9",X"3A",X"63",X"4C",X"57",X"1E",X"06",X"CD",X"F8",X"2B",X"D0",X"3A",X"F8",X"4E",
		X"CB",X"B7",X"32",X"F8",X"4E",X"C9",X"3A",X"53",X"4C",X"57",X"1E",X"05",X"CD",X"F8",X"2B",X"D0",
		X"3A",X"F8",X"4E",X"CB",X"AF",X"32",X"F8",X"4E",X"C9",X"3A",X"43",X"4C",X"57",X"1E",X"04",X"CD",
		X"F8",X"2B",X"D0",X"3A",X"F8",X"4E",X"CB",X"A7",X"32",X"F8",X"4E",X"C9",X"3A",X"33",X"4C",X"57",
		X"1E",X"03",X"CD",X"F8",X"2B",X"D0",X"3A",X"F8",X"4E",X"CB",X"9F",X"32",X"F8",X"4E",X"C9",X"3A",
		X"23",X"4C",X"57",X"1E",X"02",X"CD",X"F8",X"2B",X"D0",X"3A",X"F8",X"4E",X"CB",X"97",X"32",X"F8",
		X"4E",X"C9",X"3A",X"13",X"4C",X"57",X"1E",X"01",X"CD",X"F8",X"2B",X"D0",X"3A",X"F8",X"4E",X"CB",
		X"8F",X"32",X"F8",X"4E",X"C9",X"3A",X"03",X"4C",X"57",X"1E",X"00",X"CD",X"F8",X"2B",X"D0",X"3A",
		X"F8",X"4E",X"CB",X"87",X"32",X"F8",X"4E",X"C9",X"DD",X"7E",X"04",X"FE",X"E4",X"D2",X"21",X"2C",
		X"47",X"3E",X"E4",X"90",X"4F",X"7A",X"B9",X"38",X"0A",X"47",X"79",X"C6",X"20",X"B8",X"38",X"03",
		X"C3",X"21",X"2C",X"CD",X"F4",X"2A",X"DD",X"7E",X"13",X"E6",X"F0",X"83",X"DD",X"77",X"13",X"37",
		X"C9",X"CD",X"F4",X"2A",X"3A",X"F9",X"4E",X"E6",X"0F",X"FE",X"02",X"DA",X"3F",X"2C",X"3A",X"91",
		X"4D",X"CB",X"4F",X"CA",X"3F",X"2C",X"DD",X"7E",X"13",X"F6",X"0F",X"DD",X"77",X"13",X"C9",X"DD",
		X"7E",X"13",X"E6",X"F0",X"F6",X"0E",X"DD",X"77",X"13",X"C9",X"21",X"29",X"4D",X"22",X"89",X"4D",
		X"CD",X"8D",X"0C",X"21",X"41",X"4D",X"22",X"89",X"4D",X"CD",X"8D",X"0C",X"21",X"11",X"4D",X"22",
		X"89",X"4D",X"CD",X"8D",X"0C",X"3A",X"29",X"4F",X"A7",X"20",X"39",X"DD",X"21",X"00",X"4C",X"CD",
		X"E1",X"3B",X"DD",X"21",X"10",X"4C",X"CD",X"E1",X"3B",X"DD",X"21",X"20",X"4C",X"CD",X"E1",X"3B",
		X"DD",X"21",X"30",X"4C",X"CD",X"E1",X"3B",X"DD",X"21",X"40",X"4C",X"CD",X"E1",X"3B",X"DD",X"21",
		X"50",X"4C",X"CD",X"E1",X"3B",X"DD",X"21",X"60",X"4C",X"CD",X"E1",X"3B",X"DD",X"21",X"70",X"4C",
		X"CD",X"E1",X"3B",X"C9",X"DD",X"21",X"00",X"4C",X"CD",X"25",X"93",X"DD",X"21",X"10",X"4C",X"CD",
		X"25",X"93",X"DD",X"21",X"20",X"4C",X"CD",X"25",X"93",X"DD",X"21",X"30",X"4C",X"CD",X"25",X"93",
		X"DD",X"21",X"40",X"4C",X"CD",X"25",X"93",X"DD",X"21",X"50",X"4C",X"CD",X"25",X"93",X"DD",X"21",
		X"60",X"4C",X"CD",X"25",X"93",X"DD",X"21",X"70",X"4C",X"CD",X"25",X"93",X"C9",X"AF",X"32",X"FD",
		X"4E",X"C9",X"3A",X"FD",X"4E",X"FE",X"32",X"D4",X"DD",X"2C",X"A7",X"C2",X"35",X"2D",X"21",X"61",
		X"40",X"01",X"A0",X"00",X"7E",X"FE",X"9A",X"20",X"3C",X"09",X"7D",X"FE",X"21",X"20",X"F5",X"3A",
		X"79",X"4D",X"CB",X"7F",X"CA",X"35",X"2D",X"E6",X"CF",X"32",X"79",X"4D",X"3A",X"61",X"4D",X"CB",
		X"7F",X"CA",X"35",X"2D",X"E6",X"CF",X"32",X"61",X"4D",X"AF",X"32",X"5A",X"4D",X"32",X"72",X"4D",
		X"3A",X"53",X"4E",X"A7",X"20",X"0F",X"3A",X"7E",X"4D",X"FE",X"90",X"20",X"08",X"3A",X"66",X"4D",
		X"FE",X"90",X"CA",X"61",X"30",X"21",X"61",X"40",X"01",X"A0",X"00",X"E5",X"CD",X"A9",X"2F",X"E1",
		X"09",X"7D",X"FE",X"21",X"20",X"F5",X"3A",X"26",X"4F",X"A7",X"C0",X"DD",X"21",X"29",X"4D",X"3A",
		X"34",X"4D",X"A7",X"28",X"08",X"3A",X"2E",X"4D",X"FE",X"D4",X"D2",X"88",X"2D",X"CD",X"FA",X"2D",
		X"DD",X"21",X"41",X"4D",X"3A",X"4C",X"4D",X"A7",X"28",X"08",X"3A",X"46",X"4D",X"FE",X"D4",X"D2",
		X"88",X"2D",X"CD",X"FA",X"2D",X"21",X"29",X"4D",X"22",X"89",X"4D",X"CD",X"8D",X"0C",X"21",X"41",
		X"4D",X"22",X"89",X"4D",X"CD",X"8D",X"0C",X"C9",X"3A",X"79",X"4D",X"CB",X"7F",X"C8",X"3A",X"61",
		X"4D",X"CB",X"7F",X"C8",X"DD",X"E5",X"CD",X"93",X"31",X"DD",X"E1",X"3E",X"01",X"32",X"26",X"4F",
		X"01",X"00",X"04",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"09",X"06",X"18",X"77",X"2B",X"10",X"FC",
		X"FE",X"08",X"28",X"0A",X"F5",X"3E",X"0C",X"CD",X"CE",X"15",X"F1",X"3C",X"18",X"E2",X"21",X"59",
		X"4D",X"36",X"10",X"23",X"36",X"20",X"21",X"71",X"4D",X"36",X"10",X"23",X"36",X"20",X"3E",X"B6",
		X"32",X"61",X"4D",X"32",X"79",X"4D",X"3E",X"90",X"32",X"2F",X"4D",X"32",X"47",X"4D",X"CD",X"75",
		X"2D",X"21",X"53",X"4E",X"CB",X"C6",X"21",X"61",X"40",X"01",X"A0",X"00",X"7E",X"FE",X"9A",X"28",
		X"02",X"36",X"E1",X"09",X"7D",X"FE",X"21",X"20",X"F3",X"C9",X"DD",X"CB",X"0B",X"46",X"CA",X"AE",
		X"2E",X"DD",X"7E",X"05",X"47",X"FE",X"14",X"20",X"51",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"7E",
		X"FE",X"9A",X"28",X"11",X"FE",X"DF",X"28",X"20",X"DD",X"36",X"0B",X"00",X"DD",X"36",X"04",X"00",
		X"DD",X"36",X"05",X"F0",X"C9",X"3A",X"FC",X"4E",X"A7",X"28",X"F1",X"3D",X"32",X"FC",X"4E",X"DD",
		X"36",X"05",X"15",X"36",X"DF",X"C3",X"4C",X"2E",X"78",X"C6",X"08",X"47",X"23",X"7E",X"FE",X"DF",
		X"28",X"F6",X"2D",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"DD",X"70",X"05",X"DD",X"36",X"06",X"B8",
		X"3A",X"FB",X"4E",X"DD",X"77",X"01",X"DD",X"36",X"0B",X"01",X"DD",X"7E",X"08",X"A7",X"28",X"3B",
		X"3A",X"FE",X"4E",X"FE",X"01",X"20",X"12",X"DD",X"7E",X"06",X"FE",X"BC",X"28",X"07",X"DD",X"36",
		X"06",X"BC",X"C3",X"79",X"2E",X"DD",X"36",X"06",X"B8",X"DD",X"7E",X"05",X"D6",X"0C",X"32",X"F2",
		X"4C",X"DD",X"46",X"04",X"3E",X"F3",X"90",X"32",X"F3",X"4C",X"CD",X"D0",X"0D",X"1A",X"FE",X"DF",
		X"C8",X"3E",X"DF",X"12",X"DD",X"35",X"08",X"DD",X"34",X"09",X"C9",X"DD",X"6E",X"09",X"DD",X"66",
		X"0A",X"36",X"E0",X"DD",X"36",X"01",X"00",X"DD",X"36",X"06",X"90",X"C3",X"18",X"2E",X"DD",X"E5",
		X"DD",X"21",X"29",X"4D",X"FD",X"21",X"41",X"4D",X"2A",X"8E",X"4D",X"7E",X"E6",X"07",X"3D",X"28",
		X"3F",X"FE",X"02",X"28",X"73",X"DA",X"70",X"2F",X"DD",X"CB",X"0B",X"46",X"20",X"14",X"DD",X"36",
		X"04",X"73",X"DD",X"36",X"05",X"14",X"DD",X"36",X"08",X"06",X"DD",X"36",X"09",X"41",X"DD",X"36",
		X"0A",X"42",X"FD",X"CB",X"0B",X"46",X"C2",X"A4",X"2F",X"FD",X"36",X"04",X"9B",X"FD",X"36",X"05",
		X"14",X"FD",X"36",X"08",X"04",X"FD",X"36",X"09",X"A1",X"FD",X"36",X"0A",X"41",X"C3",X"A4",X"2F",
		X"DD",X"CB",X"0B",X"46",X"20",X"14",X"DD",X"36",X"04",X"23",X"DD",X"36",X"05",X"14",X"DD",X"36",
		X"08",X"0A",X"DD",X"36",X"09",X"81",X"DD",X"36",X"0A",X"43",X"FD",X"CB",X"0B",X"46",X"C2",X"A4",
		X"2F",X"FD",X"36",X"04",X"9B",X"FD",X"36",X"05",X"14",X"FD",X"36",X"08",X"03",X"FD",X"36",X"09",
		X"A1",X"FD",X"36",X"0A",X"41",X"C3",X"A4",X"2F",X"DD",X"CB",X"0B",X"46",X"20",X"14",X"DD",X"36",
		X"04",X"4B",X"DD",X"36",X"05",X"14",X"DD",X"36",X"08",X"08",X"DD",X"36",X"09",X"E1",X"DD",X"36",
		X"0A",X"42",X"FD",X"CB",X"0B",X"46",X"C2",X"A4",X"2F",X"FD",X"36",X"04",X"C3",X"FD",X"36",X"05",
		X"14",X"FD",X"36",X"08",X"05",X"FD",X"36",X"09",X"01",X"FD",X"36",X"0A",X"41",X"C3",X"A4",X"2F",
		X"DD",X"CB",X"0B",X"46",X"20",X"14",X"DD",X"36",X"04",X"73",X"DD",X"36",X"05",X"14",X"DD",X"36",
		X"08",X"03",X"DD",X"36",X"09",X"41",X"DD",X"36",X"0A",X"42",X"FD",X"CB",X"0B",X"46",X"20",X"14",
		X"FD",X"36",X"04",X"EB",X"FD",X"36",X"05",X"14",X"FD",X"36",X"08",X"07",X"FD",X"36",X"09",X"61",
		X"FD",X"36",X"0A",X"40",X"DD",X"E1",X"C3",X"01",X"2E",X"7E",X"FE",X"9A",X"C8",X"FE",X"DF",X"C8",
		X"FE",X"AD",X"38",X"1B",X"23",X"7E",X"FE",X"E0",X"28",X"12",X"FE",X"AA",X"38",X"0E",X"FE",X"AD",
		X"30",X"F2",X"FE",X"AC",X"28",X"03",X"3C",X"77",X"C9",X"36",X"9A",X"2B",X"36",X"AA",X"C9",X"36",
		X"9A",X"C9",X"3A",X"21",X"4F",X"A7",X"20",X"53",X"DD",X"7E",X"08",X"47",X"E6",X"30",X"FE",X"10",
		X"CA",X"DA",X"31",X"DA",X"D1",X"35",X"CB",X"78",X"CA",X"71",X"36",X"CD",X"41",X"26",X"D2",X"CA",
		X"35",X"DD",X"36",X"01",X"00",X"DD",X"36",X"05",X"00",X"DD",X"36",X"06",X"90",X"DD",X"36",X"08",
		X"C6",X"DD",X"36",X"0D",X"90",X"3A",X"22",X"4F",X"A7",X"3A",X"91",X"4D",X"20",X"0C",X"CB",X"4F",
		X"28",X"14",X"CB",X"AF",X"32",X"91",X"4D",X"C3",X"D1",X"35",X"CB",X"6F",X"28",X"08",X"CB",X"8F",
		X"32",X"91",X"4D",X"C3",X"D1",X"35",X"3E",X"01",X"32",X"21",X"4F",X"3A",X"61",X"4D",X"CB",X"7F",
		X"CA",X"71",X"36",X"3A",X"79",X"4D",X"CB",X"7F",X"CA",X"71",X"36",X"3A",X"3C",X"4D",X"CB",X"7F",
		X"C2",X"D1",X"35",X"3A",X"54",X"4D",X"CB",X"7F",X"C2",X"D1",X"35",X"3A",X"24",X"4D",X"CB",X"7F",
		X"C2",X"D1",X"35",X"3A",X"81",X"4C",X"A7",X"C2",X"D1",X"35",X"3A",X"90",X"4C",X"A7",X"C2",X"D1",
		X"35",X"3A",X"25",X"4F",X"A7",X"28",X"16",X"3A",X"29",X"4F",X"A7",X"20",X"10",X"21",X"61",X"40",
		X"01",X"A0",X"00",X"7E",X"FE",X"9A",X"C0",X"09",X"7D",X"FE",X"21",X"20",X"F6",X"CD",X"93",X"31",
		X"3A",X"25",X"4F",X"A7",X"C2",X"1D",X"31",X"3E",X"40",X"CD",X"CE",X"15",X"3A",X"89",X"4E",X"32",
		X"0B",X"4F",X"CB",X"4F",X"20",X"02",X"A7",X"C0",X"3E",X"90",X"32",X"FF",X"4C",X"DD",X"21",X"F9",
		X"4C",X"DD",X"36",X"04",X"1C",X"DD",X"36",X"05",X"0C",X"01",X"00",X"10",X"11",X"E4",X"FF",X"21",
		X"C0",X"43",X"2B",X"3A",X"FE",X"4C",X"C6",X"F8",X"32",X"FE",X"4C",X"7E",X"FE",X"BD",X"30",X"1B",
		X"7D",X"E6",X"0F",X"FE",X"0C",X"20",X"EB",X"7D",X"FE",X"5C",X"28",X"40",X"19",X"DD",X"36",X"05",
		X"0C",X"DD",X"7E",X"04",X"C6",X"08",X"DD",X"77",X"04",X"18",X"D7",X"3E",X"15",X"77",X"32",X"0B",
		X"4F",X"21",X"24",X"4F",X"CB",X"6E",X"E5",X"28",X"07",X"2A",X"A9",X"4D",X"09",X"22",X"A9",X"4D",
		X"E1",X"CB",X"4E",X"28",X"07",X"2A",X"AB",X"4D",X"09",X"22",X"AB",X"4D",X"3E",X"03",X"CD",X"CE",
		X"15",X"3E",X"B0",X"32",X"FF",X"4C",X"21",X"89",X"4E",X"CB",X"C6",X"C9",X"7C",X"FE",X"40",X"20",
		X"BB",X"3A",X"30",X"4D",X"32",X"27",X"4F",X"3A",X"48",X"4D",X"32",X"28",X"4F",X"21",X"91",X"4D",
		X"3A",X"21",X"4F",X"A7",X"28",X"04",X"CB",X"8E",X"CB",X"AE",X"3A",X"FD",X"4E",X"FE",X"32",X"D4",
		X"DD",X"2C",X"32",X"0A",X"4F",X"A7",X"20",X"02",X"CB",X"DE",X"F5",X"21",X"00",X"4C",X"CD",X"96",
		X"3A",X"21",X"10",X"4C",X"CD",X"96",X"3A",X"21",X"20",X"4C",X"CD",X"96",X"3A",X"21",X"30",X"4C",
		X"CD",X"96",X"3A",X"21",X"40",X"4C",X"CD",X"96",X"3A",X"21",X"50",X"4C",X"CD",X"96",X"3A",X"21",
		X"60",X"4C",X"CD",X"96",X"3A",X"21",X"70",X"4C",X"CD",X"96",X"3A",X"21",X"80",X"4C",X"CD",X"96",
		X"3A",X"21",X"90",X"4C",X"CD",X"96",X"3A",X"F1",X"32",X"FD",X"4E",X"3E",X"90",X"32",X"FF",X"4C",
		X"32",X"17",X"4D",X"32",X"2F",X"4D",X"32",X"47",X"4D",X"32",X"5F",X"4D",X"32",X"77",X"4D",X"32",
		X"0B",X"4F",X"C9",X"3A",X"6E",X"4E",X"A7",X"28",X"05",X"CB",X"CF",X"32",X"6E",X"4E",X"3A",X"BF",
		X"4E",X"A7",X"28",X"05",X"CB",X"CF",X"32",X"BF",X"4E",X"21",X"A4",X"4E",X"CB",X"CE",X"3E",X"90",
		X"32",X"FF",X"4C",X"3E",X"02",X"CD",X"CE",X"15",X"3E",X"9A",X"32",X"85",X"4C",X"32",X"95",X"4C",
		X"AF",X"32",X"84",X"4C",X"32",X"94",X"4C",X"21",X"80",X"4C",X"22",X"F4",X"4C",X"CD",X"16",X"0E",
		X"21",X"90",X"4C",X"22",X"F4",X"4C",X"CD",X"16",X"0E",X"C9",X"CD",X"B1",X"3A",X"3A",X"23",X"4F",
		X"F6",X"F8",X"D6",X"FA",X"CB",X"27",X"21",X"F1",X"31",X"CD",X"E3",X"15",X"5E",X"23",X"56",X"EB",
		X"E9",X"70",X"33",X"FD",X"32",X"36",X"33",X"27",X"32",X"AA",X"33",X"5A",X"34",X"8B",X"4C",X"49",
		X"5A",X"41",X"52",X"44",X"20",X"57",X"49",X"5A",X"41",X"52",X"44",X"2C",X"43",X"4F",X"50",X"59",
		X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"35",X"54",X"45",X"43",X"48",X"53",X"54",
		X"41",X"52",X"20",X"49",X"4E",X"43",X"2E",X"DD",X"7E",X"06",X"FE",X"78",X"38",X"07",X"16",X"8E",
		X"1E",X"7E",X"C3",X"39",X"32",X"16",X"76",X"1E",X"66",X"06",X"F8",X"0E",X"04",X"CD",X"D1",X"34",
		X"CA",X"26",X"35",X"DD",X"35",X"0A",X"C2",X"26",X"35",X"DD",X"7E",X"00",X"0E",X"18",X"16",X"14",
		X"1E",X"0C",X"FE",X"10",X"28",X"19",X"30",X"31",X"A7",X"C2",X"C4",X"32",X"DD",X"7E",X"01",X"A7",
		X"28",X"1F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"81",X"DD",X"77",X"00",X"C3",X"ED",X"32",X"DD",
		X"7E",X"01",X"A7",X"28",X"0C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"79",X"90",X"C3",X"69",
		X"32",X"DD",X"36",X"01",X"08",X"79",X"C3",X"69",X"32",X"BA",X"28",X"61",X"47",X"3A",X"23",X"4F",
		X"CB",X"5F",X"78",X"20",X"0B",X"FE",X"19",X"38",X"07",X"DD",X"36",X"00",X"18",X"C3",X"ED",X"32",
		X"3D",X"C3",X"69",X"32",X"BB",X"28",X"C2",X"47",X"3A",X"23",X"4F",X"CB",X"5F",X"78",X"20",X"0B",
		X"FE",X"08",X"30",X"07",X"DD",X"36",X"00",X"08",X"C3",X"ED",X"32",X"3C",X"C3",X"69",X"32",X"3E",
		X"18",X"C3",X"DB",X"32",X"47",X"3E",X"20",X"90",X"47",X"3A",X"23",X"4F",X"CB",X"5F",X"78",X"20",
		X"0A",X"FE",X"19",X"30",X"EA",X"FE",X"08",X"30",X"02",X"3E",X"08",X"DD",X"77",X"00",X"DD",X"7E",
		X"01",X"A7",X"CA",X"22",X"35",X"D6",X"08",X"DD",X"77",X"01",X"C3",X"22",X"35",X"DD",X"7E",X"01",
		X"FE",X"20",X"CA",X"22",X"35",X"C6",X"08",X"DD",X"77",X"01",X"C3",X"22",X"35",X"DD",X"7E",X"06",
		X"FE",X"78",X"38",X"07",X"16",X"8C",X"1E",X"7C",X"C3",X"0F",X"33",X"16",X"74",X"1E",X"64",X"06",
		X"F8",X"0E",X"02",X"CD",X"D1",X"34",X"CA",X"26",X"35",X"DD",X"35",X"0A",X"C2",X"26",X"35",X"DD",
		X"7E",X"00",X"0E",X"08",X"16",X"14",X"1E",X"0C",X"FE",X"10",X"CA",X"5C",X"32",X"30",X"95",X"A7",
		X"CA",X"6F",X"32",X"C3",X"A4",X"32",X"DD",X"7E",X"06",X"FE",X"78",X"38",X"07",X"16",X"7A",X"1E",
		X"8E",X"C3",X"48",X"33",X"16",X"62",X"1E",X"76",X"06",X"04",X"0E",X"03",X"CD",X"D1",X"34",X"CA",
		X"26",X"35",X"DD",X"35",X"0A",X"C2",X"26",X"35",X"DD",X"7E",X"00",X"0E",X"18",X"16",X"04",X"1E",
		X"1C",X"FE",X"10",X"CA",X"6F",X"32",X"D2",X"A4",X"32",X"A7",X"CA",X"5C",X"32",X"C3",X"A4",X"32",
		X"DD",X"7E",X"06",X"FE",X"78",X"38",X"07",X"16",X"78",X"1E",X"8C",X"C3",X"82",X"33",X"16",X"60",
		X"1E",X"74",X"06",X"04",X"0E",X"01",X"CD",X"D1",X"34",X"CA",X"26",X"35",X"DD",X"35",X"0A",X"C2",
		X"26",X"35",X"DD",X"7E",X"00",X"0E",X"08",X"16",X"04",X"1E",X"1C",X"FE",X"10",X"CA",X"5C",X"32",
		X"D2",X"C4",X"32",X"A7",X"CA",X"6F",X"32",X"C3",X"89",X"32",X"DD",X"7E",X"06",X"FE",X"78",X"38",
		X"13",X"CB",X"4F",X"CA",X"BD",X"33",X"16",X"7A",X"1E",X"8E",X"C3",X"D3",X"33",X"16",X"78",X"1E",
		X"8C",X"C3",X"D3",X"33",X"CB",X"4F",X"28",X"07",X"16",X"62",X"1E",X"76",X"C3",X"D3",X"33",X"16",
		X"60",X"1E",X"74",X"06",X"04",X"0E",X"05",X"CD",X"D1",X"34",X"CA",X"26",X"35",X"DD",X"35",X"0A",
		X"C2",X"26",X"35",X"DD",X"7E",X"00",X"0E",X"00",X"16",X"10",X"1E",X"00",X"FE",X"10",X"28",X"24",
		X"30",X"2C",X"A7",X"C2",X"42",X"34",X"DD",X"7E",X"01",X"FE",X"20",X"CA",X"22",X"35",X"C6",X"08",
		X"DD",X"77",X"01",X"C3",X"22",X"35",X"DD",X"7E",X"01",X"06",X"08",X"90",X"38",X"06",X"DD",X"77",
		X"01",X"C3",X"22",X"35",X"DD",X"36",X"01",X"08",X"DD",X"73",X"00",X"C3",X"22",X"35",X"FE",X"18",
		X"28",X"F2",X"DA",X"39",X"34",X"06",X"18",X"DD",X"71",X"00",X"90",X"CB",X"27",X"CB",X"27",X"CB",
		X"27",X"D6",X"08",X"DD",X"77",X"01",X"C3",X"22",X"35",X"47",X"3E",X"18",X"DD",X"72",X"00",X"C3",
		X"2A",X"34",X"FE",X"08",X"28",X"CE",X"D2",X"52",X"34",X"47",X"3E",X"08",X"DD",X"71",X"00",X"C3",
		X"2A",X"34",X"06",X"08",X"DD",X"72",X"00",X"C3",X"2A",X"34",X"DD",X"7E",X"06",X"FE",X"78",X"38",
		X"13",X"CB",X"4F",X"CA",X"6D",X"34",X"16",X"8E",X"1E",X"7E",X"C3",X"83",X"34",X"16",X"8C",X"1E",
		X"7C",X"C3",X"83",X"34",X"CB",X"4F",X"28",X"07",X"16",X"76",X"1E",X"66",X"C3",X"83",X"34",X"16",
		X"74",X"1E",X"64",X"06",X"F8",X"0E",X"06",X"CD",X"D1",X"34",X"CA",X"26",X"35",X"DD",X"35",X"0A",
		X"C2",X"26",X"35",X"DD",X"7E",X"00",X"0E",X"00",X"16",X"10",X"1E",X"10",X"FE",X"10",X"CA",X"BA",
		X"34",X"D2",X"1E",X"34",X"A7",X"20",X"9B",X"3A",X"23",X"4F",X"CB",X"5F",X"C2",X"06",X"34",X"DD",
		X"36",X"00",X"10",X"DD",X"36",X"01",X"10",X"C3",X"22",X"35",X"3A",X"23",X"4F",X"CB",X"5F",X"C2",
		X"F6",X"33",X"DD",X"7E",X"01",X"FE",X"10",X"D2",X"F6",X"33",X"DD",X"36",X"01",X"10",X"C3",X"22",
		X"35",X"DD",X"7E",X"08",X"E6",X"0F",X"B9",X"CA",X"07",X"35",X"21",X"6E",X"4E",X"CB",X"41",X"28",
		X"0B",X"3A",X"53",X"4E",X"A7",X"20",X"0B",X"CB",X"C6",X"C3",X"F2",X"34",X"7E",X"A7",X"28",X"02",
		X"CB",X"CE",X"DD",X"7E",X"08",X"E6",X"F0",X"81",X"DD",X"77",X"08",X"DD",X"72",X"06",X"DD",X"36",
		X"09",X"01",X"DD",X"36",X"0A",X"01",X"C9",X"DD",X"35",X"09",X"C2",X"20",X"35",X"DD",X"36",X"09",
		X"05",X"DD",X"7E",X"06",X"BB",X"28",X"05",X"80",X"DD",X"77",X"06",X"C9",X"DD",X"72",X"06",X"C9",
		X"AF",X"C9",X"DD",X"36",X"0A",X"02",X"DD",X"46",X"04",X"3E",X"F7",X"90",X"32",X"F3",X"4C",X"DD",
		X"7E",X"05",X"D6",X"08",X"32",X"F2",X"4C",X"CD",X"D0",X"0D",X"EB",X"3A",X"25",X"4F",X"A7",X"20",
		X"76",X"7E",X"FE",X"AA",X"DA",X"B7",X"35",X"FE",X"AD",X"DA",X"88",X"35",X"FE",X"D1",X"D2",X"B7",
		X"35",X"FE",X"CD",X"D2",X"94",X"35",X"DD",X"7E",X"06",X"FE",X"78",X"D2",X"B7",X"35",X"E6",X"03",
		X"C6",X"7C",X"DD",X"77",X"06",X"3A",X"29",X"4F",X"A7",X"20",X"14",X"DD",X"7E",X"04",X"D6",X"07",
		X"6F",X"DD",X"7E",X"05",X"C6",X"08",X"67",X"06",X"01",X"CD",X"D3",X"38",X"C3",X"B7",X"35",X"36",
		X"9A",X"21",X"FD",X"4E",X"35",X"C3",X"B7",X"35",X"3A",X"29",X"4F",X"A7",X"28",X"06",X"3A",X"FD",
		X"4E",X"A7",X"28",X"23",X"DD",X"36",X"00",X"10",X"DD",X"7E",X"08",X"E6",X"C0",X"F6",X"26",X"DD",
		X"77",X"08",X"DD",X"7E",X"04",X"DD",X"77",X"0B",X"DD",X"7E",X"05",X"DD",X"77",X"0C",X"DD",X"36",
		X"0D",X"98",X"21",X"53",X"4E",X"CB",X"C6",X"DD",X"CB",X"08",X"7E",X"CA",X"71",X"36",X"3A",X"23",
		X"4F",X"E6",X"10",X"CA",X"05",X"36",X"DD",X"CB",X"08",X"F6",X"DD",X"22",X"89",X"4D",X"CD",X"8D",
		X"0C",X"3A",X"FE",X"4E",X"FE",X"01",X"C0",X"DD",X"7E",X"0D",X"FE",X"90",X"C8",X"FE",X"94",X"28",
		X"18",X"FE",X"A0",X"CA",X"FE",X"35",X"D2",X"EF",X"35",X"C6",X"04",X"DD",X"77",X"0D",X"C9",X"3A",
		X"01",X"4F",X"FE",X"08",X"D8",X"DD",X"36",X"17",X"90",X"DD",X"36",X"0D",X"90",X"C9",X"DD",X"7E",
		X"17",X"DD",X"77",X"0D",X"C9",X"DD",X"CB",X"08",X"76",X"CA",X"CA",X"35",X"DD",X"CB",X"08",X"B6",
		X"DD",X"36",X"16",X"00",X"DD",X"CB",X"08",X"BE",X"DD",X"36",X"11",X"00",X"3A",X"1D",X"4E",X"A7",
		X"20",X"05",X"21",X"38",X"4E",X"CB",X"C6",X"DD",X"CB",X"06",X"4E",X"CA",X"3A",X"36",X"DD",X"CB",
		X"16",X"FE",X"DD",X"7E",X"04",X"D6",X"10",X"C3",X"42",X"36",X"DD",X"CB",X"16",X"BE",X"DD",X"7E",
		X"04",X"3C",X"DD",X"77",X"12",X"47",X"3E",X"F0",X"90",X"32",X"F3",X"4C",X"DD",X"7E",X"05",X"C6",
		X"06",X"DD",X"77",X"13",X"D6",X"10",X"32",X"F2",X"4C",X"CD",X"D0",X"0D",X"DD",X"73",X"14",X"DD",
		X"72",X"15",X"3A",X"A0",X"4C",X"C6",X"83",X"DD",X"77",X"10",X"EB",X"01",X"00",X"00",X"C3",X"D1",
		X"36",X"DD",X"7E",X"10",X"FE",X"9A",X"C2",X"C0",X"36",X"01",X"20",X"00",X"DD",X"7E",X"11",X"3D",
		X"FA",X"AC",X"36",X"DD",X"77",X"11",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"DD",X"CB",X"16",X"7E",
		X"20",X"16",X"37",X"3F",X"ED",X"42",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"36",X"9A",X"DD",X"CB",
		X"11",X"46",X"C2",X"79",X"36",X"C3",X"CA",X"35",X"09",X"C3",X"96",X"36",X"DD",X"7E",X"16",X"E6",
		X"0F",X"28",X"06",X"DD",X"35",X"16",X"C3",X"18",X"36",X"DD",X"CB",X"08",X"FE",X"C3",X"CA",X"35",
		X"DD",X"7E",X"11",X"FE",X"06",X"CA",X"80",X"37",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"01",X"20",
		X"00",X"DD",X"CB",X"16",X"7E",X"20",X"09",X"37",X"3F",X"ED",X"42",X"0E",X"08",X"C3",X"E3",X"36",
		X"09",X"0E",X"F8",X"DD",X"7E",X"12",X"FE",X"11",X"DA",X"80",X"37",X"FE",X"F1",X"D2",X"80",X"37",
		X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"3E",X"10",X"85",X"5F",
		X"54",X"3A",X"3C",X"4D",X"E6",X"70",X"FE",X"40",X"30",X"10",X"2A",X"2D",X"4D",X"7B",X"95",X"FE",
		X"11",X"30",X"07",X"7A",X"94",X"FE",X"11",X"DA",X"AD",X"37",X"3A",X"54",X"4D",X"E6",X"70",X"FE",
		X"40",X"30",X"10",X"2A",X"45",X"4D",X"7B",X"95",X"FE",X"11",X"30",X"07",X"7A",X"94",X"FE",X"11",
		X"DA",X"B6",X"37",X"3A",X"24",X"4D",X"E6",X"70",X"FE",X"40",X"30",X"0F",X"2A",X"15",X"4D",X"7B",
		X"95",X"FE",X"11",X"30",X"06",X"7A",X"94",X"FE",X"11",X"38",X"74",X"DD",X"6E",X"0E",X"DD",X"66",
		X"0F",X"7E",X"FE",X"9A",X"CA",X"37",X"38",X"E5",X"47",X"21",X"53",X"4E",X"7E",X"A7",X"20",X"07",
		X"CB",X"C6",X"3E",X"0D",X"32",X"09",X"4F",X"78",X"E1",X"FE",X"E0",X"CA",X"55",X"38",X"FE",X"AD",
		X"D2",X"5F",X"38",X"FE",X"AA",X"D2",X"80",X"38",X"FE",X"8B",X"D2",X"B5",X"38",X"C3",X"5F",X"38",
		X"DD",X"6E",X"14",X"DD",X"66",X"15",X"DD",X"75",X"0E",X"DD",X"74",X"0F",X"DD",X"36",X"10",X"9A",
		X"01",X"00",X"00",X"C3",X"7C",X"36",X"3A",X"22",X"4F",X"A7",X"C2",X"A5",X"37",X"2A",X"A9",X"4D",
		X"19",X"22",X"A9",X"4D",X"C9",X"2A",X"AB",X"4D",X"19",X"22",X"AB",X"4D",X"C9",X"DD",X"E5",X"DD",
		X"21",X"29",X"4D",X"C3",X"CA",X"37",X"DD",X"E5",X"DD",X"21",X"41",X"4D",X"C3",X"CA",X"37",X"DD",
		X"E5",X"DD",X"21",X"11",X"4D",X"21",X"A4",X"4E",X"CB",X"C6",X"3A",X"25",X"4F",X"A7",X"C2",X"00",
		X"38",X"CD",X"F4",X"2A",X"DD",X"7E",X"13",X"E6",X"80",X"F6",X"4A",X"DD",X"77",X"13",X"DD",X"36",
		X"01",X"20",X"DD",X"36",X"00",X"10",X"21",X"53",X"4E",X"CB",X"C6",X"11",X"00",X"01",X"DD",X"E1",
		X"DD",X"36",X"17",X"B4",X"CD",X"96",X"37",X"AF",X"32",X"01",X"4F",X"3E",X"98",X"C3",X"61",X"38",
		X"DD",X"36",X"01",X"00",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"F0",X"DD",X"36",X"06",X"90",
		X"DD",X"36",X"0B",X"00",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"CD",X"26",X"38",X"DD",X"E1",X"DD",
		X"36",X"17",X"B0",X"C3",X"F4",X"37",X"36",X"AA",X"7D",X"E6",X"E0",X"3C",X"6F",X"36",X"E1",X"21",
		X"FD",X"4E",X"35",X"11",X"00",X"10",X"C9",X"DD",X"7E",X"10",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",
		X"77",X"DD",X"7E",X"12",X"81",X"DD",X"77",X"12",X"DD",X"34",X"11",X"DD",X"CB",X"11",X"46",X"C2",
		X"C8",X"36",X"C3",X"CA",X"35",X"CD",X"26",X"38",X"DD",X"36",X"17",X"B0",X"C3",X"F4",X"37",X"3E",
		X"94",X"DD",X"77",X"0D",X"3E",X"06",X"32",X"FE",X"4E",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"7C",
		X"D6",X"08",X"67",X"7D",X"C6",X"08",X"6F",X"DD",X"75",X"0B",X"DD",X"74",X"0C",X"C3",X"80",X"37",
		X"3A",X"25",X"4F",X"A7",X"C2",X"80",X"37",X"3A",X"29",X"4F",X"A7",X"C2",X"AC",X"38",X"11",X"00",
		X"25",X"CD",X"96",X"37",X"06",X"01",X"DD",X"6E",X"12",X"DD",X"66",X"13",X"CD",X"D3",X"38",X"AF",
		X"32",X"01",X"4F",X"DD",X"36",X"17",X"A8",X"3E",X"98",X"C3",X"61",X"38",X"DD",X"7E",X"10",X"77",
		X"3E",X"98",X"C3",X"61",X"38",X"11",X"00",X"20",X"CD",X"96",X"37",X"06",X"00",X"DD",X"6E",X"12",
		X"DD",X"66",X"13",X"CD",X"D3",X"38",X"AF",X"32",X"01",X"4F",X"DD",X"36",X"17",X"AC",X"3E",X"98",
		X"C3",X"61",X"38",X"7D",X"FE",X"81",X"D2",X"32",X"39",X"FE",X"79",X"38",X"43",X"7C",X"FE",X"A8",
		X"DA",X"13",X"39",X"3A",X"63",X"4C",X"FE",X"78",X"30",X"08",X"3A",X"60",X"4C",X"FE",X"02",X"D2",
		X"8C",X"39",X"3A",X"43",X"4C",X"FE",X"78",X"30",X"08",X"3A",X"40",X"4C",X"FE",X"02",X"D2",X"A9",
		X"39",X"3A",X"23",X"4C",X"FE",X"78",X"30",X"08",X"3A",X"20",X"4C",X"FE",X"02",X"D2",X"C6",X"39",
		X"C3",X"E3",X"39",X"FE",X"78",X"D2",X"F2",X"38",X"FE",X"50",X"D2",X"01",X"39",X"C3",X"E3",X"39",
		X"7C",X"FE",X"A8",X"30",X"67",X"FE",X"78",X"D2",X"A9",X"39",X"FE",X"50",X"D2",X"C6",X"39",X"C3",
		X"E3",X"39",X"FE",X"89",X"30",X"43",X"7C",X"FE",X"90",X"DA",X"6C",X"39",X"3A",X"73",X"4C",X"FE",
		X"61",X"38",X"08",X"3A",X"70",X"4C",X"FE",X"02",X"D2",X"00",X"3A",X"3A",X"53",X"4C",X"FE",X"61",
		X"38",X"08",X"3A",X"50",X"4C",X"FE",X"02",X"D2",X"1D",X"3A",X"3A",X"33",X"4C",X"FE",X"61",X"38",
		X"08",X"3A",X"30",X"4C",X"FE",X"02",X"D2",X"3A",X"3A",X"C3",X"57",X"3A",X"FE",X"70",X"D2",X"4B",
		X"39",X"FE",X"48",X"D2",X"5A",X"39",X"C3",X"57",X"3A",X"7C",X"FE",X"90",X"D2",X"00",X"3A",X"FE",
		X"70",X"D2",X"1D",X"3A",X"FE",X"48",X"D2",X"3A",X"3A",X"C3",X"57",X"3A",X"78",X"FE",X"01",X"38",
		X"0C",X"21",X"F8",X"4E",X"CB",X"76",X"20",X"0C",X"0E",X"06",X"CD",X"74",X"3A",X"21",X"60",X"4C",
		X"CD",X"96",X"3A",X"C9",X"CB",X"B6",X"C3",X"9D",X"39",X"78",X"FE",X"01",X"38",X"0C",X"21",X"F8",
		X"4E",X"CB",X"66",X"20",X"0C",X"0E",X"04",X"CD",X"74",X"3A",X"21",X"40",X"4C",X"CD",X"96",X"3A",
		X"C9",X"CB",X"A6",X"C3",X"BA",X"39",X"78",X"FE",X"01",X"38",X"0C",X"21",X"F8",X"4E",X"CB",X"56",
		X"20",X"0C",X"0E",X"02",X"CD",X"74",X"3A",X"21",X"20",X"4C",X"CD",X"96",X"3A",X"C9",X"CB",X"96",
		X"C3",X"D7",X"39",X"78",X"FE",X"01",X"38",X"0C",X"21",X"F8",X"4E",X"CB",X"46",X"20",X"0C",X"0E",
		X"00",X"CD",X"74",X"3A",X"21",X"00",X"4C",X"CD",X"96",X"3A",X"C9",X"CB",X"86",X"C3",X"F4",X"39",
		X"78",X"FE",X"01",X"38",X"0C",X"21",X"F8",X"4E",X"CB",X"7E",X"20",X"0C",X"0E",X"07",X"CD",X"74",
		X"3A",X"21",X"70",X"4C",X"CD",X"96",X"3A",X"C9",X"CB",X"BE",X"C3",X"11",X"3A",X"78",X"FE",X"01",
		X"38",X"0C",X"21",X"F8",X"4E",X"CB",X"6E",X"20",X"0C",X"0E",X"05",X"CD",X"74",X"3A",X"21",X"50",
		X"4C",X"CD",X"96",X"3A",X"C9",X"CB",X"AE",X"C3",X"2E",X"3A",X"78",X"FE",X"01",X"38",X"0C",X"21",
		X"F8",X"4E",X"CB",X"5E",X"20",X"0C",X"0E",X"03",X"CD",X"74",X"3A",X"21",X"30",X"4C",X"CD",X"96",
		X"3A",X"C9",X"CB",X"9E",X"C3",X"4B",X"3A",X"78",X"FE",X"01",X"38",X"0C",X"21",X"F8",X"4E",X"CB",
		X"4E",X"20",X"0C",X"0E",X"01",X"CD",X"74",X"3A",X"21",X"10",X"4C",X"CD",X"96",X"3A",X"C9",X"CB",
		X"8E",X"C3",X"68",X"3A",X"3E",X"02",X"32",X"FA",X"4E",X"3A",X"3C",X"4D",X"47",X"E6",X"0F",X"B9",
		X"20",X"09",X"78",X"E6",X"F0",X"F6",X"0A",X"32",X"3C",X"4D",X"C9",X"3A",X"54",X"4D",X"E6",X"F0",
		X"F6",X"0A",X"32",X"54",X"4D",X"C9",X"36",X"01",X"22",X"F4",X"4C",X"DD",X"E5",X"CD",X"16",X"0E",
		X"DD",X"E1",X"AF",X"2A",X"F4",X"4C",X"23",X"23",X"23",X"77",X"23",X"77",X"21",X"FD",X"4E",X"35",
		X"C9",X"DD",X"7E",X"05",X"FE",X"11",X"DA",X"0F",X"3B",X"FE",X"CC",X"D2",X"44",X"3B",X"DD",X"7E",
		X"04",X"FE",X"20",X"DA",X"CD",X"3A",X"FE",X"F1",X"D2",X"F9",X"3A",X"3F",X"C9",X"DD",X"7E",X"00",
		X"FE",X"11",X"38",X"F7",X"47",X"DD",X"7E",X"06",X"FE",X"60",X"DA",X"E2",X"3A",X"DD",X"36",X"04",
		X"20",X"C9",X"3E",X"20",X"90",X"DD",X"77",X"00",X"DD",X"CB",X"06",X"4E",X"CA",X"F4",X"3A",X"DD",
		X"CB",X"06",X"8E",X"C9",X"DD",X"CB",X"06",X"CE",X"C9",X"DD",X"7E",X"00",X"A7",X"C8",X"FE",X"10",
		X"D0",X"47",X"DD",X"7E",X"06",X"FE",X"60",X"DA",X"E2",X"3A",X"DD",X"36",X"04",X"F0",X"C9",X"DD",
		X"7E",X"00",X"47",X"FE",X"11",X"38",X"10",X"FE",X"18",X"CA",X"BE",X"3A",X"3F",X"D0",X"3E",X"30",
		X"90",X"DD",X"77",X"00",X"C3",X"33",X"3B",X"FE",X"08",X"CA",X"BE",X"3A",X"D0",X"3E",X"10",X"90",
		X"DD",X"77",X"00",X"DD",X"7E",X"06",X"FE",X"60",X"D8",X"DD",X"7E",X"01",X"D6",X"09",X"D8",X"3C",
		X"DD",X"77",X"01",X"C9",X"DD",X"7E",X"06",X"FE",X"78",X"DA",X"C8",X"3B",X"4F",X"CB",X"4F",X"C2",
		X"C3",X"3B",X"AF",X"DD",X"86",X"04",X"47",X"FE",X"48",X"30",X"0E",X"FE",X"31",X"38",X"69",X"FE",
		X"3D",X"21",X"80",X"4C",X"38",X"22",X"C3",X"83",X"3B",X"78",X"FE",X"C1",X"38",X"5A",X"FE",X"D8",
		X"30",X"56",X"FE",X"CD",X"21",X"90",X"4C",X"38",X"05",X"06",X"20",X"C3",X"8A",X"3B",X"06",X"28",
		X"C3",X"8A",X"3B",X"06",X"B0",X"C3",X"8A",X"3B",X"06",X"B8",X"7E",X"A7",X"20",X"3A",X"79",X"D6",
		X"18",X"DD",X"77",X"06",X"36",X"03",X"23",X"23",X"23",X"70",X"23",X"36",X"C8",X"11",X"00",X"30",
		X"CD",X"96",X"37",X"3E",X"02",X"32",X"FE",X"4E",X"32",X"01",X"4F",X"DD",X"7E",X"04",X"DD",X"77",
		X"0B",X"DD",X"7E",X"05",X"DD",X"77",X"0C",X"DD",X"36",X"0D",X"A4",X"21",X"89",X"4E",X"CB",X"C6",
		X"C3",X"C8",X"3B",X"3E",X"F8",X"C3",X"53",X"3B",X"DD",X"7E",X"00",X"47",X"FE",X"11",X"38",X"08",
		X"FE",X"18",X"CA",X"BE",X"3A",X"C3",X"1D",X"3B",X"FE",X"08",X"CA",X"BE",X"3A",X"3F",X"C3",X"2C",
		X"3B",X"DD",X"22",X"F4",X"4C",X"DD",X"7E",X"00",X"FE",X"01",X"CA",X"D2",X"3C",X"D2",X"1B",X"3C",
		X"DD",X"35",X"0D",X"C0",X"DD",X"36",X"0D",X"05",X"DD",X"7E",X"05",X"FE",X"AC",X"C2",X"08",X"3C",
		X"DD",X"36",X"05",X"AA",X"CD",X"16",X"0E",X"C9",X"FE",X"AE",X"30",X"07",X"DD",X"34",X"05",X"CD",
		X"16",X"0E",X"C9",X"DD",X"36",X"05",X"AD",X"CD",X"16",X"0E",X"C9",X"DD",X"7E",X"04",X"E6",X"07",
		X"C2",X"C4",X"3C",X"DD",X"7E",X"03",X"E6",X"07",X"C2",X"C4",X"3C",X"DD",X"35",X"0D",X"C2",X"7D",
		X"3C",X"DD",X"7E",X"05",X"FE",X"8B",X"C2",X"3D",X"3C",X"DD",X"36",X"05",X"AA",X"DD",X"36",X"0D",
		X"05",X"DD",X"36",X"00",X"00",X"CD",X"16",X"0E",X"2A",X"F4",X"4C",X"7D",X"21",X"F8",X"4E",X"FE",
		X"40",X"28",X"0F",X"D2",X"6E",X"3C",X"FE",X"20",X"28",X"0E",X"30",X"09",X"A7",X"20",X"0C",X"CB",
		X"C6",X"C9",X"CB",X"E6",X"C9",X"CB",X"DE",X"C9",X"CB",X"D6",X"C9",X"CB",X"CE",X"C9",X"FE",X"60",
		X"28",X"05",X"30",X"06",X"CB",X"EE",X"C9",X"CB",X"F6",X"C9",X"CB",X"FE",X"C9",X"DD",X"7E",X"04",
		X"47",X"DD",X"7E",X"08",X"B8",X"C2",X"C4",X"3C",X"DD",X"7E",X"03",X"47",X"DD",X"7E",X"07",X"B8",
		X"C2",X"C4",X"3C",X"DD",X"6E",X"09",X"DD",X"66",X"0A",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",
		X"77",X"01",X"23",X"7E",X"DD",X"77",X"07",X"23",X"7E",X"DD",X"77",X"08",X"23",X"7E",X"23",X"FE",
		X"01",X"C2",X"C8",X"3C",X"7E",X"DD",X"77",X"09",X"23",X"7E",X"DD",X"77",X"0A",X"2A",X"8E",X"4D",
		X"7E",X"DD",X"77",X"0D",X"CD",X"16",X"0E",X"C9",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"CD",X"16",
		X"0E",X"C9",X"2A",X"F4",X"4C",X"CB",X"65",X"28",X"42",X"21",X"1F",X"4C",X"35",X"C0",X"35",X"3A",
		X"FC",X"4E",X"A7",X"C8",X"DD",X"36",X"03",X"68",X"DD",X"36",X"04",X"D0",X"3D",X"32",X"FC",X"4E",
		X"DD",X"6E",X"0B",X"DD",X"66",X"0C",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"DD",X"36",X"0D",X"00",
		X"EB",X"2A",X"8E",X"4D",X"46",X"EB",X"3A",X"FB",X"4E",X"B8",X"DA",X"14",X"3D",X"DD",X"36",X"05",
		X"8B",X"C3",X"99",X"3C",X"DD",X"36",X"05",X"AE",X"C3",X"99",X"3C",X"21",X"0F",X"4C",X"35",X"C0",
		X"35",X"3A",X"FC",X"4E",X"A7",X"C8",X"DD",X"36",X"03",X"70",X"DD",X"36",X"04",X"D0",X"C3",X"EC",
		X"3C",X"02",X"20",X"70",X"60",X"00",X"02",X"10",X"70",X"08",X"00",X"05",X"08",X"78",X"08",X"00",
		X"05",X"08",X"C0",X"08",X"00",X"03",X"08",X"C0",X"18",X"00",X"04",X"08",X"A0",X"18",X"00",X"03",
		X"08",X"A0",X"38",X"00",X"04",X"08",X"78",X"38",X"00",X"02",X"08",X"78",X"08",X"01",X"40",X"3D",
		X"02",X"20",X"68",X"60",X"00",X"02",X"10",X"68",X"10",X"00",X"04",X"08",X"60",X"10",X"00",X"04",
		X"08",X"40",X"10",X"00",X"02",X"08",X"40",X"08",X"00",X"04",X"08",X"10",X"08",X"00",X"03",X"08",
		X"10",X"18",X"00",X"05",X"08",X"30",X"18",X"00",X"03",X"08",X"30",X"30",X"00",X"05",X"08",X"60",
		X"30",X"00",X"02",X"08",X"60",X"10",X"01",X"6F",X"3D",X"02",X"20",X"70",X"60",X"00",X"02",X"10",
		X"70",X"50",X"00",X"05",X"08",X"78",X"50",X"00",X"05",X"08",X"A8",X"50",X"00",X"03",X"08",X"A8",
		X"60",X"00",X"05",X"08",X"D0",X"60",X"00",X"02",X"08",X"D0",X"48",X"00",X"04",X"08",X"90",X"48",
		X"00",X"02",X"08",X"90",X"40",X"00",X"04",X"08",X"78",X"40",X"00",X"03",X"08",X"78",X"50",X"01",
		X"A8",X"3D",X"02",X"20",X"68",X"50",X"00",X"02",X"10",X"68",X"38",X"00",X"04",X"08",X"60",X"38",
		X"00",X"04",X"08",X"38",X"38",X"00",X"03",X"08",X"38",X"48",X"00",X"04",X"08",X"08",X"48",X"00",
		X"03",X"08",X"08",X"58",X"00",X"05",X"08",X"18",X"58",X"00",X"02",X"08",X"18",X"48",X"00",X"05",
		X"08",X"28",X"48",X"00",X"03",X"08",X"28",X"58",X"00",X"05",X"08",X"40",X"58",X"00",X"02",X"08",
		X"40",X"48",X"00",X"05",X"08",X"60",X"48",X"00",X"02",X"08",X"60",X"38",X"01",X"E1",X"3D",X"02",
		X"20",X"70",X"88",X"00",X"02",X"10",X"70",X"70",X"00",X"05",X"08",X"78",X"70",X"00",X"05",X"08",
		X"80",X"70",X"00",X"02",X"08",X"80",X"68",X"00",X"05",X"08",X"A8",X"68",X"00",X"03",X"08",X"A8",
		X"80",X"00",X"04",X"08",X"98",X"80",X"00",X"03",X"08",X"98",X"90",X"00",X"04",X"08",X"88",X"90",
		X"00",X"02",X"08",X"88",X"88",X"00",X"04",X"08",X"78",X"88",X"00",X"02",X"08",X"78",X"70",X"01",
		X"2E",X"3E",X"02",X"20",X"68",X"78",X"00",X"02",X"10",X"68",X"60",X"00",X"04",X"08",X"60",X"60",
		X"00",X"03",X"08",X"60",X"78",X"00",X"04",X"08",X"38",X"78",X"00",X"02",X"08",X"38",X"70",X"00",
		X"04",X"08",X"28",X"70",X"00",X"02",X"08",X"28",X"68",X"00",X"04",X"08",X"10",X"68",X"00",X"02",
		X"08",X"10",X"60",X"00",X"05",X"08",X"60",X"60",X"01",X"71",X"3E",X"02",X"20",X"70",X"A8",X"00",
		X"02",X"10",X"70",X"98",X"00",X"05",X"08",X"78",X"98",X"00",X"05",X"08",X"A8",X"98",X"00",X"03",
		X"08",X"A8",X"B0",X"00",X"05",X"08",X"D0",X"B0",X"00",X"02",X"08",X"D0",X"98",X"00",X"04",X"08",
		X"90",X"98",X"00",X"03",X"08",X"90",X"B0",X"00",X"04",X"08",X"78",X"B0",X"00",X"02",X"08",X"78",
		X"98",X"01",X"AA",X"3E",X"02",X"20",X"68",X"98",X"00",X"02",X"10",X"68",X"80",X"00",X"04",X"08",
		X"60",X"80",X"00",X"04",X"08",X"38",X"80",X"00",X"03",X"08",X"38",X"90",X"00",X"04",X"08",X"28",
		X"90",X"00",X"03",X"08",X"28",X"98",X"00",X"04",X"08",X"08",X"98",X"00",X"03",X"08",X"08",X"B0",
		X"00",X"05",X"08",X"60",X"B0",X"00",X"02",X"08",X"60",X"A0",X"00",X"04",X"08",X"30",X"A0",X"00",
		X"02",X"08",X"30",X"98",X"00",X"05",X"08",X"60",X"98",X"00",X"02",X"08",X"60",X"80",X"01",X"E3",
		X"3E",X"3E",X"9A",X"CD",X"45",X"15",X"3E",X"02",X"CD",X"55",X"15",X"21",X"6C",X"88",X"11",X"F9",
		X"4C",X"01",X"07",X"00",X"ED",X"B0",X"21",X"84",X"88",X"11",X"11",X"4D",X"01",X"14",X"00",X"ED",
		X"B0",X"3A",X"29",X"4D",X"21",X"84",X"88",X"11",X"29",X"4D",X"01",X"14",X"00",X"ED",X"B0",X"32",
		X"29",X"4D",X"3A",X"27",X"4F",X"32",X"29",X"4D",X"3A",X"41",X"4D",X"21",X"84",X"88",X"11",X"41",
		X"4D",X"01",X"14",X"00",X"ED",X"B0",X"32",X"41",X"4D",X"3A",X"28",X"4F",X"32",X"41",X"4D",X"21",
		X"6C",X"88",X"11",X"59",X"4D",X"01",X"18",X"00",X"ED",X"B0",X"21",X"6C",X"88",X"11",X"71",X"4D",
		X"01",X"18",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"00",X"4C",X"01",X"10",X"00",X"ED",X"B0",
		X"21",X"58",X"85",X"11",X"10",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"20",
		X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"30",X"4C",X"01",X"10",X"00",X"ED",
		X"B0",X"21",X"58",X"85",X"11",X"40",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",
		X"50",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"60",X"4C",X"01",X"10",X"00",
		X"ED",X"B0",X"21",X"58",X"85",X"11",X"70",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",
		X"11",X"80",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"90",X"4C",X"01",X"10",
		X"00",X"ED",X"B0",X"3E",X"FF",X"32",X"09",X"4F",X"3E",X"D0",X"32",X"59",X"4D",X"3E",X"09",X"32");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
