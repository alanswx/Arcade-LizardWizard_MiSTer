library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"9A",X"CD",X"45",X"15",X"3E",X"02",X"CD",X"55",X"15",X"21",X"6C",X"88",X"11",X"F9",X"4C",
		X"01",X"07",X"00",X"ED",X"B0",X"21",X"84",X"88",X"11",X"11",X"4D",X"01",X"14",X"00",X"ED",X"B0",
		X"3A",X"36",X"4D",X"21",X"84",X"88",X"11",X"29",X"4D",X"01",X"14",X"00",X"ED",X"B0",X"32",X"36",
		X"4D",X"3A",X"27",X"4F",X"32",X"30",X"4D",X"3A",X"4E",X"4D",X"21",X"84",X"88",X"11",X"41",X"4D",
		X"01",X"14",X"00",X"ED",X"B0",X"32",X"4E",X"4D",X"3A",X"28",X"4F",X"32",X"48",X"4D",X"21",X"6C",
		X"88",X"11",X"59",X"4D",X"01",X"18",X"00",X"ED",X"B0",X"21",X"6C",X"88",X"11",X"71",X"4D",X"01",
		X"18",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"00",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",
		X"58",X"85",X"11",X"10",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"20",X"4C",
		X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"30",X"4C",X"01",X"10",X"00",X"ED",X"B0",
		X"21",X"58",X"85",X"11",X"40",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"50",
		X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"60",X"4C",X"01",X"10",X"00",X"ED",
		X"B0",X"21",X"58",X"85",X"11",X"70",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",
		X"80",X"4C",X"01",X"10",X"00",X"ED",X"B0",X"21",X"58",X"85",X"11",X"90",X"4C",X"01",X"10",X"00",
		X"ED",X"B0",X"3E",X"FF",X"32",X"09",X"4F",X"3E",X"D0",X"32",X"5D",X"4D",X"3E",X"09",X"32",X"60",
		X"4D",X"3D",X"32",X"1E",X"4D",X"3E",X"14",X"32",X"00",X"4D",X"3E",X"06",X"32",X"FE",X"4E",X"3E",
		X"05",X"32",X"08",X"4F",X"AF",X"32",X"80",X"4C",X"32",X"90",X"4C",X"32",X"F8",X"4E",X"32",X"F9",
		X"4E",X"32",X"FA",X"4E",X"32",X"F9",X"4C",X"32",X"FF",X"4E",X"32",X"00",X"4F",X"32",X"0B",X"4F",
		X"32",X"21",X"4F",X"32",X"25",X"4F",X"32",X"26",X"4F",X"32",X"29",X"4F",X"32",X"2A",X"4F",X"3C",
		X"32",X"0F",X"4C",X"3A",X"91",X"4D",X"32",X"24",X"4F",X"21",X"31",X"3D",X"22",X"0B",X"4C",X"21",
		X"60",X"3D",X"22",X"1B",X"4C",X"21",X"99",X"3D",X"22",X"2B",X"4C",X"21",X"D2",X"3D",X"22",X"3B",
		X"4C",X"21",X"1F",X"3E",X"22",X"4B",X"4C",X"21",X"62",X"3E",X"22",X"5B",X"4C",X"21",X"9B",X"3E",
		X"22",X"6B",X"4C",X"21",X"D4",X"3E",X"22",X"7B",X"4C",X"C9",X"11",X"8B",X"41",X"21",X"5C",X"87",
		X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"4B",X"89",X"06",X"06",X"CD",X"06",X"89",X"CD",
		X"9C",X"89",X"CD",X"98",X"88",X"CD",X"B3",X"88",X"3E",X"0C",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",
		X"A7",X"20",X"02",X"3E",X"0A",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"3E",X"6A",X"32",X"54",X"4D",
		X"3E",X"80",X"32",X"39",X"4D",X"C9",X"11",X"8B",X"41",X"21",X"65",X"87",X"3E",X"01",X"06",X"09",
		X"CD",X"66",X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"CD",X"98",X"88",X"CD",X"E9",X"88",X"06",
		X"03",X"CD",X"B7",X"89",X"3A",X"0A",X"4F",X"A7",X"20",X"02",X"3E",X"0A",X"32",X"FD",X"4E",X"32",
		X"FC",X"4E",X"3E",X"40",X"32",X"39",X"4D",X"32",X"51",X"4D",X"C9",X"11",X"8B",X"41",X"21",X"6E",
		X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"4B",X"89",X"CD",X"73",X"89",X"06",X"06",
		X"CD",X"06",X"89",X"CD",X"9C",X"89",X"CD",X"B3",X"88",X"CD",X"CE",X"88",X"06",X"04",X"CD",X"B7",
		X"89",X"3E",X"0A",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",X"A7",X"20",X"02",X"3E",X"0E",X"32",X"FD",
		X"4E",X"32",X"FC",X"4E",X"C9",X"11",X"8B",X"41",X"21",X"77",X"87",X"3E",X"01",X"06",X"09",X"CD",
		X"66",X"16",X"11",X"51",X"41",X"21",X"45",X"88",X"3E",X"03",X"06",X"0D",X"CD",X"66",X"16",X"06",
		X"06",X"CD",X"06",X"89",X"CD",X"9C",X"89",X"3A",X"91",X"4D",X"47",X"CB",X"68",X"3E",X"0C",X"28",
		X"06",X"CB",X"48",X"28",X"02",X"3E",X"11",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",X"A7",X"20",X"02",
		X"3E",X"0F",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"3E",X"0A",X"32",X"3C",X"4D",X"32",X"54",X"4D",
		X"3E",X"10",X"32",X"29",X"4D",X"32",X"41",X"4D",X"3E",X"09",X"32",X"25",X"4F",X"32",X"30",X"4D",
		X"32",X"48",X"4D",X"21",X"A4",X"4E",X"CB",X"C6",X"11",X"40",X"40",X"21",X"F0",X"86",X"3E",X"01",
		X"06",X"1C",X"CD",X"66",X"16",X"11",X"40",X"44",X"21",X"5B",X"87",X"3E",X"01",X"06",X"1C",X"CD",
		X"7C",X"16",X"21",X"91",X"4D",X"E5",X"CB",X"6E",X"28",X"09",X"21",X"77",X"4D",X"36",X"74",X"23",
		X"23",X"CB",X"E6",X"E1",X"CB",X"4E",X"C8",X"21",X"5F",X"4D",X"36",X"74",X"23",X"23",X"CB",X"E6",
		X"C9",X"11",X"8B",X"41",X"21",X"80",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"73",
		X"89",X"CD",X"81",X"89",X"06",X"06",X"CD",X"06",X"89",X"06",X"04",X"C5",X"CD",X"9C",X"89",X"CD",
		X"98",X"88",X"CD",X"B3",X"88",X"CD",X"CE",X"88",X"CD",X"E9",X"88",X"C1",X"11",X"10",X"00",X"21",
		X"01",X"4C",X"E5",X"36",X"58",X"23",X"36",X"40",X"23",X"36",X"AC",X"23",X"36",X"01",X"E1",X"19",
		X"10",X"F0",X"11",X"20",X"00",X"21",X"23",X"42",X"CD",X"5F",X"83",X"21",X"EB",X"40",X"CD",X"5F",
		X"83",X"21",X"CC",X"42",X"CD",X"5F",X"83",X"21",X"52",X"42",X"CD",X"5F",X"83",X"21",X"F3",X"40",
		X"CD",X"5F",X"83",X"3E",X"30",X"32",X"39",X"4D",X"32",X"F7",X"4E",X"3E",X"6A",X"32",X"54",X"4D",
		X"3A",X"0A",X"4F",X"A7",X"20",X"02",X"3E",X"09",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"32",X"29",
		X"4F",X"21",X"44",X"42",X"36",X"AE",X"3D",X"C8",X"21",X"A8",X"40",X"36",X"AE",X"3D",X"C8",X"21",
		X"48",X"43",X"36",X"AE",X"3D",X"C8",X"21",X"2C",X"41",X"36",X"AE",X"3D",X"C8",X"21",X"14",X"41",
		X"36",X"AE",X"3D",X"C8",X"21",X"ED",X"42",X"36",X"AE",X"3D",X"C8",X"21",X"73",X"42",X"36",X"AE",
		X"3D",X"C8",X"21",X"72",X"43",X"36",X"AE",X"3D",X"C8",X"21",X"92",X"40",X"36",X"AE",X"C9",X"E5",
		X"36",X"D8",X"19",X"36",X"D3",X"19",X"36",X"D2",X"19",X"36",X"D1",X"E1",X"01",X"00",X"04",X"09",
		X"06",X"04",X"36",X"0F",X"19",X"10",X"FB",X"C9",X"11",X"8B",X"41",X"21",X"89",X"87",X"3E",X"01",
		X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"CD",X"B3",X"88",X"CD",X"CE",
		X"88",X"CD",X"E9",X"88",X"06",X"05",X"CD",X"B7",X"89",X"3A",X"0A",X"4F",X"A7",X"20",X"02",X"3E",
		X"18",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"3E",X"0C",X"32",X"FB",X"4E",X"3E",X"03",X"32",X"08",
		X"4F",X"C9",X"11",X"8B",X"41",X"21",X"92",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",
		X"04",X"89",X"CD",X"9C",X"89",X"3A",X"91",X"4D",X"47",X"CB",X"68",X"3E",X"0E",X"28",X"06",X"CB",
		X"48",X"28",X"02",X"3E",X"13",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",X"A7",X"C2",X"42",X"82",X"3E",
		X"14",X"C3",X"42",X"82",X"11",X"8B",X"41",X"21",X"9B",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",
		X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"CD",X"CE",X"88",X"CD",X"E9",X"88",X"AF",X"32",X"FB",
		X"4E",X"3E",X"02",X"32",X"08",X"4F",X"06",X"06",X"CD",X"B7",X"89",X"3A",X"0A",X"4F",X"A7",X"20",
		X"02",X"3E",X"12",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"C9",X"11",X"8B",X"41",X"21",X"A4",X"87",
		X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"3A",X"91",X"4D",
		X"47",X"CB",X"68",X"3E",X"10",X"28",X"9E",X"CB",X"48",X"28",X"9A",X"3E",X"13",X"C3",X"D5",X"83",
		X"11",X"8B",X"41",X"21",X"AD",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",X"89",
		X"06",X"07",X"C3",X"BB",X"82",X"11",X"8B",X"41",X"21",X"B6",X"87",X"3E",X"01",X"06",X"09",X"CD",
		X"66",X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"CD",X"98",X"88",X"CD",X"B3",X"88",X"CD",X"CE",
		X"88",X"CD",X"E9",X"88",X"3E",X"0A",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",X"A7",X"20",X"02",X"3E",
		X"18",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"C9",X"3A",X"91",X"4D",X"CB",X"47",X"28",X"18",X"11",
		X"8B",X"41",X"21",X"BF",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",X"89",X"CD",
		X"CE",X"88",X"CD",X"E9",X"88",X"18",X"05",X"3E",X"09",X"CD",X"55",X"15",X"CD",X"9C",X"89",X"CD",
		X"98",X"88",X"CD",X"B3",X"88",X"3E",X"0A",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",X"A7",X"20",X"02",
		X"3E",X"18",X"32",X"FD",X"4E",X"32",X"FC",X"4E",X"C9",X"11",X"8B",X"41",X"21",X"C8",X"87",X"3E",
		X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"3A",X"91",X"4D",X"47",
		X"CB",X"68",X"3E",X"12",X"CA",X"D5",X"83",X"CB",X"48",X"CA",X"D5",X"83",X"3E",X"15",X"C3",X"D5",
		X"83",X"11",X"8B",X"41",X"21",X"D1",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",
		X"89",X"CD",X"9C",X"89",X"CD",X"98",X"88",X"CD",X"B3",X"88",X"CD",X"CE",X"88",X"CD",X"E9",X"88",
		X"3E",X"0A",X"32",X"FB",X"4E",X"3A",X"0A",X"4F",X"A7",X"20",X"02",X"3E",X"24",X"32",X"FD",X"4E",
		X"32",X"FC",X"4E",X"C9",X"11",X"8B",X"41",X"21",X"DA",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",
		X"16",X"CD",X"04",X"89",X"CD",X"9C",X"89",X"CD",X"04",X"85",X"3E",X"02",X"32",X"08",X"4F",X"C9",
		X"11",X"8B",X"41",X"21",X"E3",X"87",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"CD",X"04",X"89",
		X"CD",X"9C",X"89",X"CD",X"04",X"85",X"C9",X"C9",X"01",X"00",X"00",X"00",X"00",X"AE",X"9A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"0A",X"0B",X"0C",X"15",X"15",X"15",X"15",X"0D",
		X"0E",X"0F",X"15",X"15",X"15",X"15",X"10",X"11",X"12",X"15",X"15",X"15",X"15",X"13",X"19",X"1A",
		X"15",X"15",X"15",X"15",X"9A",X"9A",X"9A",X"15",X"15",X"15",X"15",X"9A",X"9A",X"9A",X"15",X"15",
		X"15",X"15",X"9A",X"1B",X"1C",X"15",X"15",X"15",X"15",X"9A",X"1D",X"1E",X"15",X"15",X"15",X"15",
		X"9A",X"1F",X"20",X"15",X"15",X"15",X"15",X"9A",X"21",X"22",X"15",X"15",X"15",X"23",X"24",X"25",
		X"26",X"27",X"28",X"29",X"2A",X"2B",X"2C",X"2D",X"2E",X"2F",X"5B",X"5C",X"5D",X"5E",X"5F",X"60",
		X"61",X"62",X"63",X"9A",X"14",X"64",X"65",X"66",X"67",X"16",X"9A",X"14",X"68",X"69",X"6A",X"6B",
		X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"16",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",
		X"7B",X"7C",X"7D",X"7E",X"7F",X"80",X"0A",X"0B",X"0C",X"15",X"15",X"81",X"82",X"0D",X"0E",X"0F",
		X"15",X"15",X"15",X"15",X"10",X"11",X"12",X"15",X"15",X"15",X"15",X"13",X"19",X"1A",X"15",X"15",
		X"15",X"15",X"9A",X"9A",X"9A",X"15",X"15",X"15",X"15",X"9A",X"9A",X"9A",X"15",X"15",X"15",X"15",
		X"9A",X"1B",X"1C",X"15",X"15",X"15",X"15",X"9A",X"1D",X"1E",X"15",X"15",X"15",X"15",X"9A",X"1F",
		X"20",X"15",X"15",X"15",X"15",X"9A",X"21",X"22",X"15",X"15",X"15",X"15",X"03",X"03",X"03",X"15",
		X"15",X"15",X"15",X"03",X"03",X"03",X"15",X"15",X"15",X"15",X"03",X"03",X"03",X"15",X"15",X"15",
		X"15",X"03",X"03",X"03",X"15",X"15",X"15",X"15",X"11",X"16",X"16",X"15",X"15",X"15",X"15",X"11",
		X"16",X"16",X"15",X"15",X"15",X"15",X"09",X"03",X"03",X"15",X"15",X"15",X"15",X"09",X"03",X"03",
		X"15",X"15",X"15",X"15",X"09",X"03",X"03",X"15",X"15",X"15",X"15",X"09",X"03",X"03",X"15",X"15",
		X"15",X"0E",X"03",X"03",X"0D",X"0E",X"0E",X"0E",X"0E",X"03",X"0C",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"09",X"17",X"0F",X"0F",X"0F",X"0F",X"0F",X"09",X"17",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"10",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"10",X"03",X"0D",X"0E",X"0E",X"0E",X"0F",X"03",X"03",X"03",X"15",X"15",X"0E",
		X"0E",X"03",X"03",X"03",X"15",X"15",X"15",X"15",X"03",X"03",X"03",X"15",X"15",X"15",X"15",X"03",
		X"03",X"03",X"15",X"15",X"15",X"15",X"11",X"16",X"16",X"15",X"15",X"15",X"15",X"11",X"16",X"16",
		X"15",X"15",X"15",X"15",X"09",X"03",X"03",X"15",X"15",X"15",X"15",X"09",X"03",X"03",X"15",X"15",
		X"15",X"15",X"09",X"03",X"03",X"15",X"15",X"15",X"15",X"09",X"03",X"03",X"15",X"15",X"15",X"15",
		X"D9",X"D4",X"D3",X"D3",X"D2",X"D3",X"D3",X"D1",X"D8",X"D2",X"D2",X"D3",X"D1",X"D8",X"D3",X"D3",
		X"D2",X"D3",X"D9",X"D4",X"D3",X"D3",X"D1",X"D8",X"D1",X"D8",X"D3",X"D3",X"D7",X"D6",X"D6",X"D5",
		X"9A",X"9A",X"9A",X"D4",X"9A",X"9A",X"9A",X"D3",X"9A",X"9A",X"9A",X"D2",X"9A",X"9A",X"9A",X"D1",
		X"0F",X"0F",X"0F",X"0F",X"09",X"09",X"09",X"0F",X"09",X"09",X"09",X"0F",X"09",X"09",X"09",X"0F",
		X"09",X"09",X"09",X"0F",X"9A",X"9A",X"9A",X"D8",X"9A",X"9A",X"9A",X"D3",X"9A",X"9A",X"9A",X"D2",
		X"9A",X"9A",X"9A",X"D9",X"DC",X"DB",X"DB",X"DA",X"09",X"09",X"09",X"0F",X"09",X"09",X"09",X"0F",
		X"09",X"09",X"09",X"0F",X"09",X"09",X"09",X"0F",X"0F",X"0F",X"0F",X"0F",X"31",X"40",X"40",X"40",
		X"4C",X"45",X"56",X"45",X"4C",X"32",X"40",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"33",X"40",
		X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"34",X"40",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",
		X"35",X"40",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"36",X"40",X"40",X"40",X"4C",X"45",X"56",
		X"45",X"4C",X"37",X"40",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"38",X"40",X"40",X"40",X"4C",
		X"45",X"56",X"45",X"4C",X"39",X"40",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"30",X"31",X"40",
		X"40",X"4C",X"45",X"56",X"45",X"4C",X"31",X"31",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"32",
		X"31",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"33",X"31",X"40",X"40",X"4C",X"45",X"56",X"45",
		X"4C",X"34",X"31",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"35",X"31",X"40",X"40",X"4C",X"45",
		X"56",X"45",X"4C",X"36",X"31",X"40",X"40",X"4C",X"45",X"56",X"45",X"4C",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"18",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"1B",X"1B",X"1B",X"45",X"4C",X"50",X"4F",X"45",X"50",X"40",X"45",X"55",X"43",X"53",X"45",X"52",
		X"53",X"4B",X"43",X"4F",X"52",X"40",X"54",X"4F",X"4F",X"48",X"53",X"53",X"4C",X"4C",X"41",X"42",
		X"45",X"52",X"49",X"46",X"40",X"44",X"4E",X"41",X"53",X"4E",X"4F",X"47",X"41",X"52",X"44",X"40",
		X"44",X"49",X"4F",X"56",X"41",X"53",X"40",X"53",X"52",X"59",X"52",X"4F",X"45",X"45",X"44",X"48",
		X"54",X"59",X"54",X"41",X"50",X"40",X"52",X"53",X"45",X"43",X"40",X"52",X"40",X"54",X"4F",X"48",
		X"4F",X"46",X"43",X"4F",X"45",X"55",X"48",X"42",X"4F",X"53",X"40",X"54",X"10",X"00",X"00",X"00",
		X"40",X"C8",X"90",X"08",X"C6",X"03",X"02",X"00",X"00",X"90",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"01",X"5A",X"11",X"24",X"43",X"21",X"34",X"87",X"3E",X"04",
		X"06",X"05",X"CD",X"66",X"16",X"11",X"24",X"47",X"21",X"48",X"87",X"3E",X"04",X"06",X"05",X"CD",
		X"66",X"16",X"C9",X"11",X"44",X"40",X"21",X"0C",X"87",X"3E",X"04",X"06",X"05",X"CD",X"66",X"16",
		X"11",X"44",X"44",X"21",X"20",X"87",X"3E",X"04",X"06",X"05",X"CD",X"66",X"16",X"C9",X"11",X"2E",
		X"43",X"21",X"34",X"87",X"3E",X"04",X"06",X"05",X"CD",X"66",X"16",X"11",X"2E",X"47",X"21",X"48",
		X"87",X"3E",X"04",X"06",X"05",X"CD",X"66",X"16",X"C9",X"11",X"4E",X"40",X"21",X"0C",X"87",X"3E",
		X"04",X"06",X"05",X"CD",X"66",X"16",X"11",X"4E",X"44",X"21",X"20",X"87",X"3E",X"04",X"06",X"05",
		X"CD",X"66",X"16",X"C9",X"06",X"03",X"C5",X"11",X"8B",X"45",X"21",X"EC",X"87",X"3E",X"01",X"06",
		X"09",X"CD",X"66",X"16",X"3E",X"0A",X"CD",X"CE",X"15",X"11",X"8B",X"45",X"21",X"01",X"88",X"3E",
		X"01",X"06",X"09",X"CD",X"66",X"16",X"3E",X"0A",X"CD",X"CE",X"15",X"11",X"8B",X"45",X"21",X"0A",
		X"88",X"3E",X"01",X"06",X"09",X"CD",X"66",X"16",X"3E",X"0A",X"CD",X"CE",X"15",X"C1",X"10",X"C6",
		X"3E",X"9A",X"CD",X"45",X"15",X"3E",X"09",X"CD",X"55",X"15",X"C9",X"11",X"73",X"41",X"21",X"20",
		X"88",X"3E",X"01",X"06",X"0B",X"CD",X"66",X"16",X"11",X"55",X"41",X"21",X"2B",X"88",X"3E",X"01",
		X"06",X"0D",X"CD",X"66",X"16",X"11",X"59",X"41",X"21",X"38",X"88",X"3E",X"01",X"06",X"0D",X"CD",
		X"66",X"16",X"C9",X"11",X"4F",X"41",X"21",X"13",X"88",X"3E",X"01",X"06",X"0D",X"CD",X"66",X"16",
		X"C9",X"11",X"56",X"41",X"21",X"38",X"88",X"3E",X"01",X"06",X"0D",X"CD",X"66",X"16",X"11",X"58",
		X"41",X"21",X"2B",X"88",X"3E",X"01",X"06",X"0D",X"CD",X"66",X"16",X"C9",X"11",X"59",X"40",X"21",
		X"68",X"85",X"3E",X"07",X"06",X"1C",X"CD",X"66",X"16",X"11",X"59",X"44",X"21",X"2C",X"86",X"3E",
		X"07",X"06",X"1C",X"CD",X"66",X"16",X"C9",X"3A",X"36",X"4D",X"B8",X"30",X"04",X"78",X"32",X"36",
		X"4D",X"3A",X"4E",X"4D",X"B8",X"D0",X"78",X"32",X"4E",X"4D",X"C9",X"32",X"C9",X"C9",X"3E",X"E2",
		X"01",X"16",X"08",X"18",X"05",X"3E",X"40",X"01",X"00",X"00",X"32",X"FE",X"4E",X"21",X"40",X"40",
		X"AF",X"32",X"03",X"4F",X"11",X"BF",X"43",X"7D",X"FE",X"ED",X"28",X"0B",X"FE",X"C0",X"20",X"0C",
		X"7C",X"FE",X"43",X"28",X"5B",X"18",X"05",X"7C",X"FE",X"41",X"28",X"4C",X"C5",X"46",X"3A",X"FE",
		X"4E",X"B8",X"C1",X"28",X"4B",X"CD",X"62",X"8A",X"3A",X"02",X"4F",X"3C",X"32",X"02",X"4F",X"E6",
		X"07",X"20",X"09",X"C5",X"E5",X"3E",X"01",X"CD",X"CE",X"15",X"E1",X"C1",X"3A",X"03",X"4F",X"FE",
		X"02",X"28",X"15",X"30",X"1F",X"A7",X"28",X"04",X"23",X"1B",X"18",X"BB",X"C5",X"01",X"20",X"00",
		X"09",X"EB",X"ED",X"42",X"C1",X"EB",X"18",X"AF",X"C5",X"EB",X"01",X"20",X"00",X"09",X"EB",X"ED",
		X"42",X"C1",X"18",X"A3",X"2B",X"13",X"18",X"9F",X"3A",X"FE",X"4E",X"FE",X"40",X"20",X"86",X"C9",
		X"3A",X"03",X"4F",X"3C",X"E6",X"03",X"32",X"03",X"4F",X"2A",X"04",X"4F",X"ED",X"5B",X"06",X"4F",
		X"18",X"A6",X"77",X"22",X"04",X"4F",X"F5",X"78",X"CD",X"75",X"8A",X"F1",X"77",X"22",X"06",X"4F",
		X"79",X"CD",X"75",X"8A",X"C9",X"C5",X"01",X"00",X"04",X"09",X"77",X"ED",X"42",X"C1",X"EB",X"C9",
		X"C9",X"21",X"CC",X"8B",X"22",X"8E",X"4D",X"3E",X"12",X"32",X"0A",X"4F",X"3E",X"04",X"32",X"36",
		X"4D",X"32",X"4E",X"4D",X"3E",X"07",X"32",X"27",X"4F",X"32",X"28",X"4F",X"C9",X"3E",X"FF",X"32",
		X"F5",X"4D",X"C9",X"AF",X"32",X"36",X"4D",X"32",X"4E",X"4D",X"32",X"FF",X"4E",X"32",X"00",X"4F",
		X"32",X"0A",X"4F",X"CD",X"55",X"15",X"3E",X"15",X"CD",X"45",X"15",X"3E",X"07",X"32",X"27",X"4F",
		X"32",X"28",X"4F",X"3E",X"D0",X"32",X"F7",X"4E",X"C9",X"11",X"47",X"40",X"21",X"83",X"92",X"3E",
		X"02",X"06",X"1B",X"CD",X"66",X"16",X"11",X"47",X"44",X"21",X"84",X"8B",X"3E",X"02",X"06",X"1B",
		X"CD",X"7C",X"16",X"11",X"4B",X"40",X"21",X"B9",X"92",X"3E",X"04",X"06",X"1B",X"CD",X"66",X"16",
		X"11",X"4B",X"44",X"21",X"85",X"8B",X"3E",X"04",X"06",X"1B",X"CD",X"7C",X"16",X"11",X"51",X"40",
		X"21",X"18",X"8B",X"3E",X"04",X"06",X"1B",X"CD",X"66",X"16",X"11",X"51",X"44",X"21",X"86",X"8B",
		X"3E",X"04",X"06",X"1B",X"CD",X"7C",X"16",X"C9",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"40",X"54",X"4C",X"40",X"48",X"45",X"4C",X"55",X"43",X"4E",X"49",X"4F",X"41",X"41",X"57",X"59",
		X"45",X"4C",X"40",X"40",X"40",X"50",X"53",X"54",X"45",X"40",X"44",X"53",X"53",X"4F",X"52",X"4E",
		X"49",X"54",X"41",X"49",X"52",X"40",X"5A",X"41",X"41",X"44",X"49",X"47",X"40",X"45",X"4C",X"41",
		X"45",X"55",X"40",X"40",X"4C",X"43",X"45",X"4D",X"50",X"53",X"48",X"45",X"4F",X"45",X"54",X"48",
		X"45",X"52",X"40",X"54",X"50",X"40",X"52",X"40",X"40",X"45",X"4F",X"45",X"45",X"42",X"40",X"56",
		X"48",X"40",X"53",X"41",X"54",X"54",X"55",X"4C",X"40",X"53",X"46",X"53",X"53",X"55",X"59",X"4E",
		X"41",X"4D",X"5A",X"45",X"1A",X"02",X"18",X"00",X"00",X"15",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"45",X"00",X"00",X"00",X"60",X"00",X"00",X"50",X"12",X"00",X"00",X"00",X"25",X"00",X"00",
		X"50",X"37",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"40",X"00",X"00",X"50",X"07",X"00",X"00",X"00",X"15",X"00",X"00",
		X"50",X"22",X"00",X"00",X"00",X"30",X"00",X"05",X"04",X"03",X"02",X"01",X"02",X"03",X"04",X"09",
		X"0A",X"0B",X"0C",X"FF",X"4D",X"49",X"43",X"50",X"42",X"03",X"4C",X"4C",X"44",X"60",X"17",X"03",
		X"4C",X"52",X"53",X"20",X"85",X"02",X"42",X"49",X"4C",X"90",X"76",X"02",X"41",X"4E",X"47",X"50",
		X"31",X"02",X"42",X"55",X"42",X"90",X"10",X"02",X"44",X"4F",X"43",X"00",X"05",X"02",X"46",X"4C",
		X"4F",X"60",X"01",X"02",X"4A",X"52",X"46",X"80",X"98",X"01",X"52",X"41",X"59",X"40",X"86",X"01",
		X"1B",X"18",X"1A",X"00",X"C7",X"FA",X"00",X"A0",X"FE",X"00",X"9B",X"EE",X"00",X"8B",X"FE",X"00",
		X"6B",X"EE",X"00",X"5D",X"FC",X"00",X"17",X"EB",X"00",X"15",X"FF",X"00",X"33",X"EB",X"00",X"81",
		X"FB",X"00",X"A3",X"EB",X"01",X"D2",X"FA",X"00",X"C5",X"FE",X"00",X"8C",X"FD",X"00",X"80",X"FF",
		X"00",X"CA",X"FC",X"00",X"C1",X"EC",X"00",X"A9",X"FE",X"00",X"6E",X"EE",X"00",X"26",X"FC",X"00",
		X"1C",X"EC",X"00",X"19",X"FD",X"00",X"6B",X"FF",X"00",X"9A",X"FB",X"00",X"CA",X"FA",X"00",X"91",
		X"EE",X"00",X"2E",X"FD",X"00",X"50",X"FF",X"00",X"C9",X"FB",X"00",X"15",X"0B",X"1D",X"4E",X"0B",
		X"38",X"4E",X"0C",X"02",X"01",X"43",X"00",X"02",X"08",X"05",X"04",X"01",X"54",X"00",X"05",X"04",
		X"01",X"32",X"00",X"05",X"04",X"01",X"85",X"00",X"05",X"04",X"01",X"A7",X"00",X"05",X"04",X"01",
		X"64",X"00",X"05",X"04",X"01",X"0B",X"01",X"05",X"04",X"09",X"0B",X"02",X"4E",X"0B",X"38",X"4E",
		X"01",X"F0",X"00",X"0C",X"02",X"06",X"02",X"0F",X"05",X"03",X"02",X"00",X"05",X"03",X"07",X"0F",
		X"09",X"0C",X"07",X"02",X"0F",X"01",X"00",X"01",X"06",X"06",X"05",X"01",X"03",X"F0",X"FF",X"07",
		X"06",X"03",X"50",X"00",X"04",X"FE",X"07",X"06",X"09",X"0B",X"6E",X"4E",X"0B",X"89",X"4E",X"0C",
		X"02",X"01",X"40",X"00",X"02",X"0F",X"06",X"05",X"01",X"03",X"F0",X"FF",X"07",X"02",X"05",X"03",
		X"01",X"70",X"00",X"06",X"05",X"01",X"03",X"F0",X"FF",X"07",X"06",X"02",X"08",X"01",X"00",X"0A",
		X"0C",X"06",X"06",X"05",X"02",X"03",X"E0",X"FF",X"07",X"38",X"09",X"0C",X"06",X"01",X"60",X"00",
		X"02",X"0C",X"06",X"06",X"06",X"05",X"01",X"03",X"10",X"00",X"07",X"06",X"03",X"A0",X"FF",X"07",
		X"02",X"04",X"FF",X"07",X"0B",X"09",X"0B",X"53",X"4E",X"0B",X"6E",X"4E",X"0C",X"06",X"02",X"0F",
		X"01",X"00",X"00",X"06",X"03",X"1A",X"00",X"05",X"01",X"07",X"0E",X"09",X"0B",X"BF",X"4E",X"0C",
		X"02",X"06",X"01",X"58",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"58",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"02",X"01",X"05",X"0C",X"01",X"43",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"07",X"02",X"01",X"58",X"00",X"02",
		X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"43",X"00",X"02",X"08",X"06",X"05",X"02",
		X"04",X"FF",X"07",X"05",X"01",X"58",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",
		X"01",X"64",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"06",X"01",X"69",X"00",
		X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"69",X"00",X"02",X"08",X"06",X"05",
		X"02",X"04",X"FF",X"07",X"05",X"02",X"01",X"05",X"0C",X"01",X"4F",X"00",X"02",X"08",X"06",X"05",
		X"02",X"04",X"FF",X"07",X"05",X"07",X"02",X"01",X"69",X"00",X"02",X"08",X"06",X"05",X"02",X"04",
		X"FF",X"07",X"05",X"01",X"4F",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",
		X"69",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"76",X"00",X"02",X"08",
		X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"06",X"01",X"7D",X"00",X"02",X"08",X"06",X"05",X"02",
		X"04",X"FF",X"07",X"05",X"01",X"7D",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",
		X"02",X"01",X"05",X"0C",X"01",X"5E",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",
		X"07",X"02",X"01",X"7D",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"5E",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"76",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"5E",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"05",X"06",X"01",X"70",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",
		X"70",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"02",X"01",X"05",X"0C",X"01",
		X"54",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"07",X"02",X"01",X"70",X"00",
		X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"54",X"00",X"02",X"08",X"06",X"05",
		X"02",X"04",X"FF",X"07",X"05",X"01",X"69",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",
		X"05",X"01",X"54",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"06",X"01",X"64",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"64",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"05",X"02",X"01",X"05",X"0C",X"01",X"4B",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"05",X"07",X"02",X"01",X"64",X"00",X"02",X"08",X"06",X"05",X"02",
		X"04",X"FF",X"07",X"05",X"01",X"4B",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",
		X"01",X"5E",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"01",X"4B",X"00",X"02",
		X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"05",X"08",X"31",X"8D",X"09",X"0B",X"A4",X"4E",X"0C",
		X"02",X"02",X"0F",X"01",X"00",X"01",X"06",X"03",X"18",X"00",X"05",X"01",X"07",X"0C",X"05",X"02",
		X"08",X"03",X"8F",X"09",X"0C",X"02",X"01",X"58",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"58",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"70",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"70",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"85",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"85",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"95",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"95",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"76",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"76",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"95",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"95",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"B1",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"B1",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"C7",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"C7",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"85",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"85",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"A7",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"A7",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"C7",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"C7",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"E0",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"C7",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"0B",X"01",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",
		X"07",X"03",X"01",X"C7",X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"E0",
		X"00",X"02",X"08",X"06",X"05",X"02",X"04",X"FF",X"07",X"03",X"01",X"B1",X"00",X"02",X"08",X"06",
		X"05",X"02",X"04",X"FF",X"07",X"06",X"05",X"0C",X"09",X"3E",X"88",X"32",X"0C",X"4F",X"3E",X"9A",
		X"CD",X"45",X"15",X"3E",X"08",X"CD",X"55",X"15",X"CD",X"9C",X"89",X"CD",X"98",X"88",X"CD",X"B3",
		X"88",X"11",X"24",X"41",X"21",X"75",X"92",X"3E",X"01",X"06",X"0E",X"CD",X"66",X"16",X"11",X"24",
		X"45",X"21",X"EC",X"87",X"3E",X"01",X"06",X"0E",X"CD",X"66",X"16",X"3E",X"3C",X"CD",X"CE",X"15",
		X"11",X"09",X"43",X"21",X"47",X"92",X"3E",X"04",X"06",X"04",X"CD",X"66",X"16",X"11",X"0F",X"43",
		X"21",X"57",X"92",X"3E",X"04",X"06",X"04",X"CD",X"66",X"16",X"11",X"89",X"40",X"21",X"F7",X"91",
		X"3E",X"04",X"06",X"14",X"CD",X"66",X"16",X"11",X"8F",X"40",X"21",X"F7",X"91",X"3E",X"04",X"06",
		X"14",X"CD",X"66",X"16",X"11",X"37",X"41",X"21",X"67",X"92",X"3E",X"01",X"06",X"0E",X"CD",X"66",
		X"16",X"11",X"37",X"45",X"21",X"EC",X"87",X"3E",X"01",X"06",X"0E",X"CD",X"66",X"16",X"3A",X"90",
		X"4D",X"CB",X"6F",X"C0",X"21",X"10",X"4F",X"34",X"21",X"0D",X"4F",X"3A",X"0C",X"43",X"FE",X"AB",
		X"38",X"0C",X"28",X"14",X"36",X"AA",X"23",X"36",X"AB",X"23",X"36",X"AC",X"18",X"12",X"36",X"AB",
		X"23",X"36",X"AC",X"23",X"36",X"AA",X"18",X"08",X"36",X"AC",X"23",X"36",X"AA",X"23",X"36",X"AB",
		X"11",X"09",X"43",X"21",X"47",X"92",X"CD",X"EC",X"91",X"11",X"8F",X"41",X"21",X"17",X"92",X"CD",
		X"94",X"91",X"11",X"0F",X"43",X"21",X"57",X"92",X"CD",X"94",X"91",X"11",X"89",X"40",X"21",X"F7",
		X"91",X"CD",X"EC",X"91",X"11",X"0F",X"41",X"21",X"07",X"92",X"CD",X"94",X"91",X"11",X"89",X"42",
		X"21",X"37",X"92",X"CD",X"94",X"91",X"11",X"8F",X"40",X"21",X"F7",X"91",X"CD",X"EC",X"91",X"11",
		X"09",X"41",X"21",X"07",X"92",X"CD",X"94",X"91",X"11",X"0F",X"42",X"21",X"27",X"92",X"CD",X"94",
		X"91",X"11",X"89",X"41",X"21",X"17",X"92",X"CD",X"EC",X"91",X"11",X"8F",X"42",X"21",X"37",X"92",
		X"CD",X"94",X"91",X"11",X"09",X"42",X"21",X"27",X"92",X"CD",X"94",X"91",X"21",X"0C",X"4F",X"34",
		X"C2",X"EE",X"90",X"C9",X"D5",X"11",X"11",X"4F",X"D5",X"06",X"10",X"7E",X"FE",X"9A",X"28",X"3E",
		X"FE",X"3F",X"30",X"17",X"4F",X"3A",X"10",X"4F",X"CB",X"47",X"79",X"28",X"31",X"FE",X"3C",X"28",
		X"19",X"38",X"13",X"FE",X"3E",X"28",X"1B",X"3E",X"3E",X"18",X"23",X"FE",X"AB",X"38",X"17",X"28",
		X"1A",X"3A",X"0F",X"4F",X"18",X"18",X"3E",X"3C",X"18",X"14",X"3E",X"3B",X"18",X"10",X"3E",X"3E",
		X"18",X"0C",X"3E",X"3D",X"18",X"08",X"3A",X"0D",X"4F",X"18",X"03",X"3A",X"0E",X"4F",X"12",X"13",
		X"23",X"10",X"B8",X"E1",X"D1",X"3E",X"04",X"47",X"CD",X"66",X"16",X"C9",X"3E",X"01",X"E5",X"CD",
		X"CE",X"15",X"E1",X"CD",X"94",X"91",X"C9",X"9A",X"AA",X"AB",X"9A",X"AC",X"9A",X"9A",X"AA",X"AB",
		X"AC",X"AA",X"AB",X"9A",X"9A",X"9A",X"9A",X"9A",X"AA",X"9A",X"AC",X"AB",X"9A",X"AC",X"9A",X"AA",
		X"AC",X"AB",X"AA",X"9A",X"9A",X"9A",X"9A",X"9A",X"AA",X"AC",X"AB",X"AB",X"9A",X"AA",X"9A",X"9A",
		X"AC",X"AB",X"AA",X"9A",X"9A",X"9A",X"9A",X"AA",X"3E",X"9A",X"AB",X"AC",X"3C",X"3D",X"AA",X"AB",
		X"9A",X"3B",X"AC",X"9A",X"9A",X"9A",X"9A",X"AA",X"9A",X"9A",X"AA",X"AC",X"AB",X"AA",X"AB",X"AB",
		X"9A",X"9A",X"AC",X"9A",X"9A",X"9A",X"9A",X"9A",X"9A",X"9A",X"AA",X"9A",X"9A",X"9A",X"AB",X"9A",
		X"9A",X"9A",X"AC",X"AA",X"AC",X"AA",X"AB",X"AA",X"AC",X"AB",X"3E",X"9A",X"9A",X"3D",X"3C",X"9A",
		X"9A",X"3B",X"3D",X"AB",X"AC",X"AA",X"3B",X"52",X"41",X"54",X"53",X"48",X"43",X"45",X"54",X"40",
		X"35",X"38",X"39",X"31",X"18",X"53",X"54",X"4E",X"45",X"53",X"45",X"52",X"50",X"40",X"40",X"4E",
		X"4E",X"55",X"53",X"54",X"40",X"48",X"40",X"47",X"40",X"55",X"40",X"41",X"53",X"43",X"55",X"40",
		X"46",X"45",X"59",X"4C",X"5A",X"50",X"40",X"4F",X"54",X"45",X"45",X"50",X"4E",X"40",X"41",X"45",
		X"4C",X"48",X"50",X"54",X"40",X"40",X"45",X"45",X"48",X"45",X"54",X"52",X"40",X"46",X"4E",X"40",
		X"49",X"50",X"48",X"4C",X"54",X"45",X"49",X"48",X"57",X"40",X"4C",X"40",X"40",X"40",X"4C",X"40",
		X"40",X"40",X"49",X"40",X"45",X"45",X"57",X"45",X"52",X"48",X"40",X"42",X"49",X"54",X"59",X"40",
		X"46",X"40",X"45",X"44",X"40",X"54",X"48",X"4E",X"52",X"4F",X"54",X"41",X"4F",X"4F",X"40",X"40",
		X"46",X"48",X"52",X"53",X"40",X"53",X"4F",X"45",X"53",X"40",X"40",X"4D",X"44",X"54",X"53",X"41",
		X"52",X"53",X"4B",X"4C",X"41",X"55",X"43",X"46",X"5A",X"4D",X"4F",X"40",X"49",X"40",X"52",X"4F",
		X"4C",X"55",X"40",X"54",X"40",X"4F",X"47",X"4E",X"59",X"59",X"4E",X"49",X"42",X"40",X"49",X"40",
		X"40",X"54",X"54",X"54",X"4E",X"53",X"50",X"53",X"45",X"52",X"55",X"52",X"54",X"49",X"52",X"55",
		X"41",X"46",X"45",X"42",X"45",X"DD",X"22",X"F4",X"4C",X"DD",X"CB",X"04",X"46",X"C8",X"DD",X"6E",
		X"01",X"DD",X"66",X"02",X"7E",X"FE",X"8B",X"30",X"04",X"FE",X"83",X"30",X"1C",X"3A",X"FE",X"4E",
		X"FE",X"03",X"28",X"03",X"FE",X"06",X"C0",X"DD",X"34",X"03",X"DD",X"7E",X"03",X"FE",X"AC",X"DD",
		X"6E",X"01",X"DD",X"66",X"02",X"30",X"11",X"77",X"C9",X"36",X"9A",X"DD",X"36",X"01",X"58",X"DD",
		X"36",X"02",X"40",X"DD",X"36",X"03",X"AC",X"C9",X"36",X"9A",X"23",X"7D",X"E6",X"1F",X"FE",X"1A",
		X"30",X"5C",X"7E",X"FE",X"9A",X"20",X"11",X"DD",X"36",X"00",X"01",X"36",X"AA",X"DD",X"75",X"01",
		X"DD",X"74",X"02",X"DD",X"36",X"03",X"AA",X"C9",X"FE",X"D1",X"38",X"42",X"FE",X"DD",X"30",X"3E",
		X"DD",X"7E",X"00",X"FE",X"01",X"28",X"18",X"38",X"0B",X"01",X"DF",X"FF",X"09",X"DD",X"36",X"00",
		X"02",X"C3",X"7B",X"93",X"01",X"1F",X"00",X"09",X"DD",X"36",X"00",X"00",X"C3",X"7B",X"93",X"7D",
		X"E6",X"1F",X"FE",X"07",X"28",X"10",X"FE",X"11",X"28",X"0C",X"EB",X"2A",X"8E",X"4D",X"CB",X"46",
		X"EB",X"28",X"E1",X"C3",X"99",X"93",X"7C",X"FE",X"42",X"38",X"D9",X"C3",X"99",X"93",X"21",X"06",
		X"4C",X"35",X"C0",X"36",X"0C",X"2A",X"8E",X"4D",X"7E",X"FE",X"09",X"28",X"20",X"38",X"4E",X"FE",
		X"0B",X"28",X"32",X"30",X"52",X"3A",X"05",X"4C",X"FE",X"04",X"C8",X"DD",X"36",X"01",X"A0",X"DD",
		X"36",X"02",X"41",X"DD",X"36",X"03",X"A9",X"3E",X"04",X"32",X"05",X"4C",X"C9",X"3A",X"05",X"4C",
		X"FE",X"06",X"C8",X"DD",X"36",X"01",X"60",X"DD",X"36",X"02",X"40",X"DD",X"36",X"03",X"A9",X"3E",
		X"06",X"32",X"05",X"4C",X"C9",X"3A",X"05",X"4C",X"FE",X"02",X"C8",X"DD",X"36",X"01",X"E0",X"DD",
		X"36",X"02",X"42",X"DD",X"36",X"03",X"A9",X"3E",X"02",X"32",X"05",X"4C",X"C9",X"FE",X"02",X"28",
		X"1E",X"38",X"34",X"FE",X"03",X"20",X"DE",X"3A",X"05",X"4C",X"FE",X"05",X"C8",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"41",X"DD",X"36",X"03",X"A9",X"3E",X"05",X"32",X"05",X"4C",X"C9",X"3A",
		X"05",X"4C",X"FE",X"03",X"C8",X"DD",X"36",X"01",X"40",X"DD",X"36",X"02",X"42",X"DD",X"36",X"03",
		X"A9",X"3E",X"03",X"32",X"05",X"4C",X"C9",X"3A",X"05",X"4C",X"FE",X"01",X"C8",X"DD",X"36",X"01",
		X"80",X"DD",X"36",X"02",X"43",X"DD",X"36",X"03",X"A9",X"3E",X"01",X"32",X"05",X"4C",X"C9",X"4C",
		X"FF",X"11",X"F2",X"43",X"CD",X"ED",X"15",X"21",X"92",X"4D",X"CB",X"86",X"3E",X"01",X"CD",X"70",
		X"15",X"C9",X"D1",X"3E",X"80",X"CD",X"52",X"16",X"3E",X"20",X"CD",X"52",X"16",X"18",X"D9",X"3A",
		X"F7",X"4D",X"FE",X"00",X"CA",X"16",X"14",X"3D",X"32",X"F7",X"4D",X"FE",X"1A",X"28",X"14",X"3E",
		X"1B",X"2A",X"F9",X"4D",X"77",X"3E",X"20",X"CD",X"E3",X"15",X"22",X"F9",X"4D",X"3E",X"1A",X"77",
		X"C3",X"16",X"14",X"3D",X"32",X"F7",X"4D",X"3E",X"1B",X"2A",X"F9",X"4D",X"2B",X"77",X"23",X"77",
		X"23",X"77",X"2B",X"3E",X"40",X"18",X"E0",X"3A",X"F7",X"4D",X"FE",X"1B",X"CA",X"16",X"14",X"3C",
		X"32",X"F7",X"4D",X"FE",X"1A",X"28",X"14",X"3E",X"1B",X"2A",X"F9",X"4D",X"77",X"3E",X"20",X"CD",
		X"48",X"16",X"22",X"F9",X"4D",X"3E",X"1A",X"77",X"C3",X"16",X"14",X"3C",X"32",X"F7",X"4D",X"3E",
		X"1B",X"2A",X"F9",X"4D",X"77",X"3E",X"40",X"CD",X"48",X"16",X"22",X"F9",X"4D",X"3E",X"1A",X"2B",
		X"77",X"23",X"77",X"23",X"77",X"C3",X"16",X"14",X"3E",X"08",X"CD",X"CE",X"15",X"32",X"C0",X"50",
		X"06",X"14",X"CD",X"90",X"15",X"DA",X"4E",X"14",X"C3",X"FF",X"13",X"3A",X"F5",X"4D",X"21",X"92",
		X"4D",X"CB",X"66",X"28",X"03",X"3A",X"F6",X"4D",X"CB",X"67",X"32",X"C0",X"50",X"28",X"EC",X"18",
		X"DC",X"02",X"1B",X"18",X"1A",X"21",X"40",X"40",X"11",X"41",X"40",X"01",X"7F",X"03",X"77",X"ED",
		X"B0",X"32",X"C0",X"50",X"C9",X"21",X"40",X"44",X"11",X"41",X"44",X"01",X"7F",X"03",X"77",X"ED",
		X"B0",X"32",X"C0",X"50",X"C9",X"3E",X"02",X"CD",X"55",X"15",X"3E",X"40",X"CD",X"45",X"15",X"C9",
		X"47",X"AF",X"32",X"99",X"4D",X"32",X"9B",X"4D",X"3A",X"9B",X"4D",X"B8",X"C8",X"21",X"90",X"4D",
		X"CB",X"6E",X"C0",X"32",X"C0",X"50",X"18",X"F0",X"E5",X"21",X"20",X"00",X"19",X"EB",X"E1",X"C9",
		X"3A",X"92",X"4D",X"CB",X"47",X"28",X"0D",X"3A",X"9C",X"4D",X"47",X"3A",X"9B",X"4D",X"B8",X"30",
		X"19",X"37",X"3F",X"C9",X"78",X"32",X"9C",X"4D",X"3A",X"92",X"4D",X"CB",X"C7",X"32",X"92",X"4D",
		X"AF",X"32",X"9B",X"4D",X"32",X"99",X"4D",X"37",X"3F",X"C9",X"3A",X"92",X"4D",X"CB",X"87",X"32",
		X"92",X"4D",X"37",X"C9",X"21",X"90",X"4D",X"CB",X"FE",X"CB",X"7E",X"C8",X"18",X"FB",X"47",X"AF",
		X"32",X"9A",X"4D",X"3A",X"9A",X"4D",X"B8",X"C8",X"21",X"90",X"4D",X"CB",X"6E",X"C0",X"32",X"C0",
		X"50",X"18",X"F0",X"85",X"6F",X"D0",X"24",X"C9",X"83",X"5F",X"D0",X"14",X"C9",X"3E",X"03",X"F5",
		X"7E",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"47",X"3A",X"91",X"4D",X"CB",
		X"77",X"28",X"22",X"78",X"12",X"1B",X"7E",X"E6",X"0F",X"47",X"3A",X"91",X"4D",X"CB",X"77",X"32",
		X"91",X"4D",X"28",X"20",X"78",X"12",X"2B",X"1B",X"F1",X"3D",X"20",X"D3",X"3A",X"91",X"4D",X"CB",
		X"B7",X"32",X"91",X"4D",X"C9",X"78",X"FE",X"00",X"28",X"DB",X"3A",X"91",X"4D",X"CB",X"F7",X"32",
		X"91",X"4D",X"18",X"CF",X"78",X"FE",X"00",X"28",X"DD",X"3A",X"91",X"4D",X"CB",X"F7",X"32",X"91",
		X"4D",X"18",X"D1",X"81",X"4F",X"D0",X"04",X"C9",X"D5",X"16",X"00",X"5F",X"37",X"3F",X"ED",X"52",
		X"D1",X"C9",X"E5",X"EB",X"16",X"00",X"5F",X"37",X"3F",X"ED",X"52",X"EB",X"E1",X"C9",X"CD",X"5B",
		X"1A",X"DD",X"CB",X"00",X"D6",X"C9",X"32",X"F8",X"4C",X"D5",X"3A",X"F8",X"4C",X"4F",X"ED",X"A0",
		X"79",X"FE",X"00",X"20",X"F9",X"D1",X"CD",X"88",X"15",X"10",X"EE",X"C9",X"32",X"F8",X"4C",X"D5",
		X"3A",X"F8",X"4C",X"4F",X"ED",X"A0",X"2B",X"79",X"FE",X"00",X"20",X"F8",X"D1",X"CD",X"88",X"15",
		X"10",X"ED",X"C9",X"DD",X"7E",X"05",X"FD",X"96",X"05",X"B8",X"DA",X"E5",X"16",X"57",X"3E",X"FF",
		X"90",X"47",X"7A",X"B8",X"D2",X"E5",X"16",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"B9",X"DA",X"0F",
		X"17",X"57",X"3E",X"FF",X"91",X"4F",X"7A",X"B9",X"D2",X"0F",X"17",X"FD",X"7E",X"05",X"DD",X"BE",
		X"05",X"D2",X"24",X"17",X"FD",X"7E",X"04",X"DD",X"BE",X"04",X"D2",X"2C",X"17",X"3A",X"FF",X"4D",
		X"21",X"DD",X"16",X"CB",X"27",X"CD",X"E3",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"A9",X"17",X"82",
		X"17",X"34",X"17",X"5B",X"17",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"B9",X"38",X"18",X"57",X"3E",
		X"FF",X"91",X"4F",X"7A",X"B9",X"30",X"0F",X"DD",X"7E",X"04",X"FD",X"BE",X"04",X"38",X"0A",X"DD",
		X"36",X"00",X"18",X"3E",X"02",X"C9",X"3E",X"01",X"C9",X"DD",X"36",X"00",X"08",X"18",X"F4",X"DD",
		X"7E",X"05",X"FD",X"BE",X"05",X"38",X"07",X"DD",X"36",X"00",X"00",X"3E",X"03",X"C9",X"DD",X"36",
		X"00",X"10",X"18",X"F7",X"21",X"FF",X"4D",X"CB",X"C6",X"C3",X"C4",X"16",X"21",X"FF",X"4D",X"CB",
		X"CE",X"C3",X"CD",X"16",X"FD",X"7E",X"04",X"DD",X"96",X"04",X"47",X"DD",X"7E",X"05",X"FD",X"96",
		X"05",X"B8",X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",X"02",X"C3",X"CD",X"17",X"DD",X"36",X"00",
		X"04",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"06",X"C3",X"CD",X"17",X"FD",X"7E",X"04",X"DD",X"96",
		X"04",X"47",X"FD",X"7E",X"05",X"DD",X"96",X"05",X"B8",X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",
		X"0E",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"0C",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"0A",X"C3",
		X"CD",X"17",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"47",X"FD",X"7E",X"05",X"DD",X"96",X"05",X"B8",
		X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",X"12",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"14",X"C3",
		X"CD",X"17",X"DD",X"36",X"00",X"16",X"C3",X"CD",X"17",X"DD",X"7E",X"04",X"FD",X"96",X"04",X"47",
		X"DD",X"7E",X"05",X"FD",X"96",X"05",X"B8",X"28",X"09",X"38",X"0E",X"DD",X"36",X"00",X"1E",X"C3",
		X"CD",X"17",X"DD",X"36",X"00",X"1C",X"C3",X"CD",X"17",X"DD",X"36",X"00",X"1A",X"AF",X"32",X"FF",
		X"4D",X"C9",X"2A",X"FD",X"4D",X"E5",X"21",X"13",X"8C",X"7D",X"E1",X"BD",X"CC",X"0F",X"18",X"7E",
		X"FE",X"00",X"CA",X"F5",X"17",X"23",X"46",X"3A",X"75",X"4D",X"B8",X"CA",X"05",X"18",X"2B",X"22",
		X"FD",X"4D",X"C3",X"0E",X"18",X"23",X"46",X"3A",X"76",X"4D",X"B8",X"CA",X"05",X"18",X"2B",X"22",
		X"FD",X"4D",X"C3",X"0E",X"18",X"23",X"7E",X"32",X"F5",X"4D",X"23",X"22",X"FD",X"4D",X"C9",X"3E",
		X"FF",X"32",X"F5",X"4D",X"C9",X"3A",X"00",X"50",X"E6",X"0F",X"47",X"3A",X"40",X"50",X"E6",X"F0",
		X"B0",X"32",X"F5",X"4D",X"C9",X"3A",X"40",X"50",X"47",X"E6",X"0F",X"CB",X"78",X"28",X"02",X"CB",
		X"E7",X"32",X"F6",X"4D",X"C9",X"DD",X"21",X"02",X"4E",X"DD",X"CB",X"00",X"46",X"C4",X"5E",X"16",
		X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"51",X"50",X"CD",X"5E",X"19",
		X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"1D",X"4E",X"DD",X"CB",X"00",X"46",X"C4",X"5E",
		X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"51",X"50",X"CD",X"5E",
		X"19",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"38",X"4E",X"DD",X"CB",X"00",X"46",X"C4",
		X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"51",X"50",X"CD",
		X"5E",X"19",X"DD",X"7E",X"06",X"32",X"45",X"50",X"DD",X"21",X"53",X"4E",X"DD",X"CB",X"00",X"46",
		X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"56",X"50",
		X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"6E",X"4E",X"DD",X"CB",X"00",
		X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",X"56",
		X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"89",X"4E",X"DD",X"CB",
		X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",X"21",
		X"56",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4A",X"50",X"DD",X"21",X"A4",X"4E",X"DD",
		X"CB",X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",X"FD",
		X"21",X"5B",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4F",X"50",X"DD",X"21",X"BF",X"4E",
		X"DD",X"CB",X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"28",X"10",X"CD",X"87",X"19",
		X"FD",X"21",X"5B",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4F",X"50",X"DD",X"21",X"DA",
		X"4E",X"DD",X"CB",X"00",X"46",X"C4",X"5E",X"16",X"DD",X"CB",X"00",X"56",X"C8",X"CD",X"87",X"19",
		X"FD",X"21",X"5B",X"50",X"CD",X"5E",X"19",X"DD",X"7E",X"06",X"32",X"4F",X"50",X"C9",X"DD",X"7E",
		X"03",X"FD",X"77",X"00",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FD",X"77",X"01",X"DD",
		X"7E",X"04",X"FD",X"77",X"02",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"FD",X"77",X"03",
		X"DD",X"7E",X"05",X"FD",X"77",X"04",X"C9",X"DD",X"CB",X"00",X"4E",X"C2",X"5B",X"1A",X"DD",X"6E",
		X"01",X"DD",X"66",X"02",X"7E",X"CB",X"27",X"11",X"A5",X"19",X"CD",X"E8",X"15",X"23",X"E5",X"1A",
		X"6F",X"13",X"1A",X"67",X"E9",X"BF",X"19",X"C3",X"19",X"D1",X"19",X"DA",X"19",X"F0",X"19",X"FD",
		X"19",X"17",X"1A",X"30",X"1A",X"52",X"1A",X"5A",X"1A",X"79",X"1A",X"85",X"1A",X"91",X"1A",X"E1",
		X"C3",X"94",X"19",X"E1",X"7E",X"DD",X"77",X"03",X"23",X"7E",X"23",X"DD",X"77",X"04",X"C3",X"94",
		X"19",X"E1",X"7E",X"DD",X"77",X"05",X"23",X"C3",X"94",X"19",X"E1",X"7E",X"DD",X"46",X"03",X"80",
		X"DD",X"77",X"03",X"23",X"7E",X"23",X"DD",X"46",X"04",X"88",X"DD",X"77",X"04",X"C3",X"94",X"19",
		X"E1",X"7E",X"DD",X"46",X"05",X"80",X"DD",X"77",X"05",X"23",X"C3",X"94",X"19",X"E1",X"DD",X"7E",
		X"07",X"BE",X"30",X"0B",X"DD",X"34",X"07",X"2B",X"DD",X"75",X"01",X"DD",X"74",X"02",X"C9",X"DD",
		X"36",X"07",X"00",X"23",X"C3",X"94",X"19",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"D1",X"D5",X"2B",
		X"72",X"2B",X"73",X"2B",X"36",X"00",X"DD",X"75",X"08",X"DD",X"74",X"09",X"E1",X"C3",X"94",X"19",
		X"D1",X"1A",X"DD",X"6E",X"08",X"DD",X"66",X"09",X"BE",X"28",X"09",X"34",X"23",X"5E",X"23",X"56",
		X"EB",X"C3",X"94",X"19",X"23",X"23",X"23",X"DD",X"75",X"08",X"DD",X"74",X"09",X"13",X"EB",X"C3",
		X"94",X"19",X"E1",X"5E",X"23",X"56",X"EB",X"C3",X"94",X"19",X"E1",X"DD",X"E5",X"DD",X"E5",X"E1",
		X"D1",X"13",X"36",X"00",X"01",X"18",X"00",X"ED",X"B0",X"1A",X"DD",X"77",X"01",X"13",X"1A",X"DD",
		X"77",X"02",X"DD",X"75",X"08",X"DD",X"74",X"09",X"C9",X"E1",X"DD",X"75",X"01",X"DD",X"74",X"02",
		X"DD",X"36",X"00",X"00",X"C9",X"E1",X"5E",X"23",X"56",X"EB",X"36",X"06",X"13",X"EB",X"C3",X"94",
		X"19",X"E1",X"7E",X"DD",X"77",X"06",X"23",X"C3",X"94",X"19",X"32",X"40",X"52",X"45",X"59",X"41",
		X"4C",X"50",X"40",X"45",X"52",X"4F",X"43",X"53",X"50",X"4F",X"54",X"40",X"31",X"40",X"52",X"45",
		X"59",X"41",X"4C",X"50",X"54",X"49",X"44",X"45",X"52",X"43",X"59",X"41",X"4C",X"50",X"45",X"45",
		X"52",X"46",X"40",X"4E",X"49",X"4F",X"43",X"40",X"54",X"52",X"45",X"53",X"4E",X"49",X"52",X"45",
		X"59",X"41",X"4C",X"50",X"40",X"45",X"4E",X"4F",X"40",X"54",X"43",X"45",X"4C",X"45",X"53",X"52",
		X"4F",X"53",X"52",X"45",X"59",X"41",X"4C",X"50",X"40",X"4F",X"57",X"54",X"40",X"52",X"4F",X"40",
		X"45",X"4E",X"4F",X"40",X"54",X"43",X"45",X"4C",X"45",X"53",X"50",X"55",X"40",X"45",X"4E",X"4F",
		X"40",X"52",X"45",X"59",X"41",X"4C",X"50",X"50",X"55",X"40",X"4F",X"57",X"54",X"40",X"52",X"45",
		X"59",X"41",X"4C",X"50",X"52",X"45",X"56",X"4F",X"40",X"45",X"4D",X"41",X"47",X"59",X"52",X"44",
		X"52",X"41",X"5A",X"49",X"57",X"40",X"46",X"4F",X"40",X"4C",X"4C",X"41",X"48",X"45",X"48",X"54",
		X"40",X"4E",X"49",X"40",X"53",X"49",X"40",X"45",X"52",X"4F",X"43",X"53",X"40",X"52",X"55",X"4F",
		X"59",X"4E",X"45",X"54",X"40",X"50",X"4F",X"54",X"54",X"43",X"45",X"4C",X"45",X"53",X"40",X"4F",
		X"54",X"40",X"4B",X"43",X"49",X"54",X"53",X"59",X"4F",X"4A",X"40",X"45",X"53",X"55",X"4E",X"4F",
		X"54",X"54",X"55",X"42",X"40",X"45",X"52",X"49",X"46",X"40",X"44",X"4E",X"41",X"40",X"52",X"45",
		X"54",X"54",X"45",X"4C",X"54",X"4E",X"49",X"52",X"50",X"40",X"4F",X"54",X"45",X"4E",X"44",X"4D",
		X"41",X"4C",X"53",X"53",X"4E",X"4F",X"49",X"54",X"43",X"55",X"52",X"54",X"53",X"4E",X"49",X"40",
		X"59",X"41",X"4C",X"50",X"40",X"31",X"40",X"53",X"4E",X"49",X"4F",X"43",X"40",X"32",X"53",X"59",
		X"41",X"4C",X"50",X"40",X"32",X"40",X"40",X"4E",X"49",X"4F",X"43",X"40",X"31",X"40",X"59",X"41",
		X"4C",X"50",X"40",X"31",X"40",X"40",X"4E",X"49",X"4F",X"43",X"40",X"31",X"53",X"54",X"4E",X"49",
		X"4F",X"50",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"59",X"52",X"45",X"56",X"45",X"40",
		X"53",X"55",X"4E",X"4F",X"42",X"30",X"30",X"30",X"30",X"35",X"31",X"30",X"30",X"30",X"35",X"32",
		X"31",X"30",X"30",X"30",X"30",X"30",X"31",X"40",X"30",X"30",X"30",X"35",X"37",X"53",X"43",X"49",
		X"54",X"53",X"4F",X"4E",X"47",X"41",X"49",X"44",X"4E",X"4F",X"49",X"54",X"49",X"44",X"4E",X"4F",
		X"43",X"40",X"40",X"4E",X"4F",X"49",X"54",X"41",X"43",X"4F",X"4C",X"40",X"40",X"4D",X"4F",X"52",
		X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"44",X"37",X"40",X"40",X"40",
		X"40",X"40",X"40",X"31",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"46",
		X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"32",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"48",X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"33",X"44",X"4F",X"4F",X"47",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4A",X"37",X"40",X"40",X"40",X"40",X"40",X"40",X"34",
		X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"48",X"34",X"40",X"40",X"40",
		X"40",X"40",X"40",X"31",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4C",
		X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"32",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",
		X"40",X"40",X"40",X"4A",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"33",X"44",X"4F",X"4F",X"47",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4D",X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"34",
		X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4B",X"34",X"40",X"40",X"40",
		X"40",X"40",X"40",X"35",X"44",X"4F",X"4F",X"47",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"4E",
		X"34",X"40",X"40",X"40",X"40",X"40",X"40",X"36",X"44",X"41",X"42",X"40",X"4E",X"4F",X"49",X"54",
		X"49",X"44",X"4E",X"4F",X"43",X"40",X"40",X"4E",X"4F",X"49",X"54",X"41",X"43",X"4F",X"4C",X"40",
		X"40",X"4D",X"41",X"52",X"4E",X"45",X"4D",X"40",X"41",X"52",X"54",X"58",X"45",X"40",X"32",X"40",
		X"52",X"4F",X"46",X"06",X"03",X"1A",X"BE",X"38",X"08",X"20",X"0E",X"2B",X"1B",X"10",X"F6",X"18",
		X"06",X"CD",X"1E",X"1D",X"37",X"3F",X"C9",X"37",X"C9",X"CD",X"1E",X"1D",X"37",X"C9",X"78",X"FE",
		X"00",X"C8",X"2B",X"1B",X"3D",X"20",X"FB",X"C9",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",
		X"08",X"09",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"4A",X"4B",X"4C",X"4D",X"4E",
		X"4F",X"50",X"51",X"52",X"53",X"54",X"55",X"56",X"57",X"58",X"59",X"5A",X"5A",X"59",X"58",X"57",
		X"56",X"55",X"54",X"53",X"52",X"51",X"50",X"4F",X"4E",X"4D",X"4C",X"4B",X"4A",X"49",X"48",X"47",
		X"46",X"45",X"44",X"43",X"42",X"41",X"00",X"01",X"04",X"02",X"94",X"42",X"95",X"42",X"96",X"42",
		X"97",X"42",X"98",X"42",X"99",X"42",X"9A",X"42",X"9B",X"42",X"9C",X"42",X"9D",X"42",X"03",X"02",
		X"01",X"00",X"00",X"80",X"60",X"40",X"3A",X"FD",X"4E",X"A7",X"20",X"15",X"21",X"BF",X"4E",X"CB",
		X"56",X"28",X"0E",X"3A",X"2A",X"4F",X"3C",X"32",X"2A",X"4F",X"20",X"05",X"CB",X"CE",X"C3",X"11",
		X"31",X"3A",X"0B",X"4F",X"A7",X"C2",X"8C",X"30",X"21",X"09",X"4F",X"CB",X"7E",X"20",X"0E",X"35",
		X"20",X"0B",X"3A",X"53",X"4E",X"A7",X"28",X"05",X"CB",X"CF",X"32",X"53",X"4E",X"3A",X"77",X"4D",
		X"FE",X"78",X"DA",X"CA",X"1D",X"FE",X"90",X"DA",X"D7",X"1D",X"3A",X"5F",X"4D",X"FE",X"78",X"DA",
		X"0A",X"1E",X"FE",X"90",X"D2",X"0A",X"1E",X"3A",X"FE",X"4E",X"FE",X"01",X"C2",X"17",X"1E",X"3A",
		X"39",X"43",X"FE",X"E4",X"DA",X"F9",X"1D",X"3E",X"DD",X"32",X"39",X"43",X"32",X"F9",X"40",X"3C",
		X"32",X"19",X"43",X"32",X"D9",X"40",X"C3",X"17",X"1E",X"3E",X"E4",X"32",X"39",X"43",X"32",X"19",
		X"43",X"32",X"F9",X"40",X"32",X"D9",X"40",X"C3",X"17",X"1E",X"3A",X"39",X"43",X"FE",X"9A",X"CA",
		X"17",X"1E",X"3E",X"9A",X"C3",X"FB",X"1D",X"3A",X"80",X"4C",X"A7",X"CA",X"36",X"1E",X"DD",X"21",
		X"80",X"4C",X"21",X"A4",X"1E",X"3A",X"81",X"4C",X"A7",X"CA",X"58",X"1E",X"CD",X"6D",X"1E",X"DD",
		X"22",X"F4",X"4C",X"CD",X"16",X"0E",X"3A",X"90",X"4C",X"A7",X"CA",X"39",X"20",X"21",X"BC",X"1E",
		X"DD",X"21",X"90",X"4C",X"3A",X"91",X"4C",X"A7",X"CA",X"58",X"1E",X"CD",X"6D",X"1E",X"DD",X"22",
		X"F4",X"4C",X"CD",X"16",X"0E",X"C3",X"39",X"20",X"DD",X"36",X"01",X"10",X"DD",X"36",X"05",X"AE",
		X"DD",X"7E",X"09",X"CB",X"27",X"CD",X"E3",X"15",X"5E",X"23",X"56",X"EB",X"E9",X"DD",X"7E",X"04",
		X"DD",X"96",X"08",X"C0",X"DD",X"7E",X"03",X"DD",X"96",X"07",X"CA",X"8A",X"1E",X"DA",X"85",X"1E",
		X"DD",X"36",X"00",X"04",X"C9",X"DD",X"36",X"00",X"05",X"C9",X"DD",X"36",X"00",X"00",X"DD",X"36",
		X"01",X"00",X"2A",X"8E",X"4D",X"CB",X"46",X"CA",X"9F",X"1E",X"DD",X"36",X"05",X"BE",X"C9",X"DD",
		X"36",X"05",X"BD",X"C9",X"D4",X"1E",X"E3",X"1E",X"F2",X"1E",X"01",X"1F",X"10",X"1F",X"1F",X"1F",
		X"2E",X"1F",X"3D",X"1F",X"4C",X"1F",X"5B",X"1F",X"6A",X"1F",X"79",X"1F",X"88",X"1F",X"97",X"1F",
		X"A6",X"1F",X"B5",X"1F",X"C4",X"1F",X"D3",X"1F",X"E2",X"1F",X"F1",X"1F",X"00",X"20",X"0F",X"20",
		X"1E",X"20",X"2D",X"20",X"DD",X"36",X"07",X"D0",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"01",
		X"C3",X"36",X"1E",X"DD",X"36",X"07",X"98",X"DD",X"36",X"08",X"E8",X"DD",X"36",X"09",X"02",X"C3",
		X"36",X"1E",X"DD",X"36",X"07",X"C8",X"DD",X"36",X"08",X"E8",X"DD",X"36",X"09",X"03",X"C3",X"36",
		X"1E",X"DD",X"36",X"07",X"D0",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"04",X"C3",X"36",X"1E",
		X"DD",X"36",X"07",X"A0",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"05",X"C3",X"36",X"1E",X"DD",
		X"36",X"07",X"A0",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"06",X"C3",X"36",X"1E",X"DD",X"36",
		X"07",X"D8",X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"07",X"C3",X"36",X"1E",X"DD",X"36",X"07",
		X"B8",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"08",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"A8",
		X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"09",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"C8",X"DD",
		X"36",X"08",X"F0",X"DD",X"36",X"09",X"0A",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"B0",X"DD",X"36",
		X"08",X"E8",X"DD",X"36",X"09",X"0B",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"B8",X"DD",X"36",X"08",
		X"E0",X"DD",X"36",X"09",X"0B",X"C3",X"36",X"1E",X"DD",X"36",X"07",X"08",X"DD",X"36",X"08",X"F8",
		X"DD",X"36",X"09",X"01",X"C3",X"39",X"20",X"DD",X"36",X"07",X"40",X"DD",X"36",X"08",X"E8",X"DD",
		X"36",X"09",X"02",X"C3",X"39",X"20",X"DD",X"36",X"07",X"10",X"DD",X"36",X"08",X"E8",X"DD",X"36",
		X"09",X"03",X"C3",X"39",X"20",X"DD",X"36",X"07",X"08",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",
		X"04",X"C3",X"39",X"20",X"DD",X"36",X"07",X"38",X"DD",X"36",X"08",X"E0",X"DD",X"36",X"09",X"05",
		X"C3",X"39",X"20",X"DD",X"36",X"07",X"38",X"DD",X"36",X"08",X"F8",X"DD",X"36",X"09",X"06",X"C3",
		X"39",X"20",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"F0",X"DD",X"36",X"09",X"07",X"C3",X"39",
		X"20",X"DD",X"36",X"07",X"20",X"DD",X"36",X"7D",X"F8",X"DD",X"36",X"09",X"08",X"C3",X"39",X"0A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
