library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"22",X"00",X"00",X"00",
		X"11",X"99",X"DD",X"DD",X"FF",X"77",X"33",X"00",X"33",X"77",X"55",X"44",X"44",X"66",X"22",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"33",X"22",X"00",X"44",X"66",X"77",X"55",X"44",X"44",X"00",X"00",
		X"44",X"FF",X"FF",X"44",X"44",X"CC",X"CC",X"00",X"00",X"77",X"77",X"66",X"33",X"11",X"00",X"00",
		X"EE",X"FF",X"11",X"11",X"11",X"33",X"22",X"00",X"00",X"55",X"55",X"55",X"55",X"77",X"77",X"00",
		X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",X"00",
		X"00",X"00",X"88",X"FF",X"77",X"00",X"00",X"00",X"66",X"77",X"55",X"44",X"44",X"66",X"66",X"00",
		X"66",X"77",X"DD",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"77",X"33",X"00",
		X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",X"00",
		X"10",X"00",X"30",X"70",X"F0",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"C3",X"E1",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",
		X"00",X"00",X"00",X"01",X"01",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"70",X"3C",X"0F",X"1F",X"3F",X"3F",X"1F",X"0F",
		X"0F",X"0F",X"8F",X"CF",X"EF",X"FF",X"FF",X"FF",X"E3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"03",X"03",X"01",X"03",X"0F",X"0F",X"0F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"0F",X"7F",X"7F",X"FF",X"3F",X"3F",X"3F",X"1F",
		X"FF",X"FF",X"FF",X"FC",X"F8",X"F8",X"F8",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"07",X"07",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"7F",X"7F",X"7F",X"7E",X"3C",X"78",X"F0",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"F0",
		X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FC",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"30",X"32",X"77",X"70",X"F0",X"F0",X"10",X"00",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"E1",X"C3",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E1",
		X"77",X"77",X"77",X"EF",X"CF",X"0F",X"8F",X"CF",X"00",X"00",X"00",X"00",X"11",X"11",X"77",X"77",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E9",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"11",X"11",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E9",X"CF",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"FC",X"F8",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"10",X"30",X"70",X"F0",X"F0",
		X"87",X"C3",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"30",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"10",X"10",X"00",X"30",X"70",X"F0",
		X"F0",X"F0",X"87",X"0F",X"87",X"87",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"E0",X"00",X"01",X"83",X"00",X"FE",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"33",X"00",X"84",X"86",X"FF",X"FF",X"FF",X"00",X"00",X"0E",X"0E",X"78",
		X"FF",X"FF",X"FF",X"CC",X"00",X"00",X"0F",X"E1",X"FF",X"FF",X"FF",X"FF",X"88",X"00",X"00",X"03",
		X"00",X"00",X"07",X"0F",X"0F",X"0E",X"00",X"F0",X"EE",X"CC",X"88",X"00",X"01",X"0F",X"0C",X"10",
		X"07",X"0F",X"69",X"F0",X"C3",X"87",X"87",X"0F",X"00",X"07",X"0F",X"3C",X"78",X"70",X"F0",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"00",X"00",X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"07",X"00",X"60",X"F0",X"F0",X"F0",X"EE",X"CC",X"CC",X"EE",X"CC",X"88",X"10",X"F0",
		X"00",X"70",X"30",X"00",X"C0",X"F0",X"F0",X"F0",X"00",X"00",X"E0",X"F0",X"30",X"30",X"30",X"10",
		X"0C",X"00",X"C1",X"C3",X"C3",X"E1",X"E1",X"F0",X"0F",X"1F",X"F0",X"F0",X"10",X"C0",X"F0",X"F0",
		X"00",X"03",X"0F",X"78",X"30",X"00",X"00",X"08",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"01",X"0F",X"88",X"00",X"00",X"00",X"10",X"10",X"D0",X"C3",X"33",X"00",X"00",
		X"FE",X"FA",X"EC",X"C0",X"00",X"00",X"00",X"00",X"80",X"30",X"C4",X"10",X"00",X"00",X"00",X"00",
		X"FC",X"F5",X"EE",X"40",X"00",X"00",X"00",X"00",X"00",X"54",X"A8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"80",X"E8",X"FE",X"F4",X"00",X"00",X"00",X"00",X"00",X"50",X"11",X"FD",
		X"00",X"00",X"00",X"00",X"60",X"F6",X"F9",X"F6",X"00",X"00",X"00",X"00",X"44",X"91",X"00",X"71",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"0F",X"0F",X"F0",X"F0",X"00",X"80",X"00",X"00",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"3C",X"F0",X"F0",X"F0",X"30",X"10",X"00",X"00",
		X"11",X"33",X"33",X"00",X"00",X"33",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",X"FF",X"FF",
		X"F0",X"70",X"70",X"30",X"30",X"30",X"10",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"FF",X"FF",X"CC",
		X"F0",X"F0",X"F0",X"C0",X"00",X"F0",X"F0",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",
		X"C0",X"F0",X"F0",X"E0",X"00",X"10",X"F0",X"87",X"1E",X"1E",X"F0",X"70",X"00",X"F0",X"F0",X"F0",
		X"00",X"30",X"F0",X"87",X"0F",X"0F",X"87",X"3C",X"00",X"00",X"30",X"70",X"30",X"10",X"F0",X"0F",
		X"00",X"00",X"00",X"F0",X"96",X"0F",X"0F",X"F0",X"00",X"00",X"F0",X"F0",X"3C",X"0F",X"E1",X"F0",
		X"84",X"07",X"F0",X"F0",X"F0",X"F0",X"70",X"30",X"98",X"00",X"30",X"70",X"70",X"70",X"00",X"CC",
		X"0F",X"00",X"0C",X"0F",X"0F",X"0F",X"87",X"F0",X"0C",X"08",X"0F",X"E1",X"C3",X"F0",X"F0",X"F0",
		X"87",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C3",X"F0",X"F0",X"70",X"F0",X"1E",X"0F",X"3C",X"F0",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"1E",
		X"00",X"0E",X"E0",X"F0",X"F0",X"F0",X"F0",X"10",X"CC",X"01",X"01",X"03",X"30",X"30",X"00",X"88",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"80",X"30",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"C3",X"F0",X"F0",X"F0",X"F0",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"3C",X"96",X"C3",X"E1",X"F0",X"F0",X"1E",X"87",X"E1",X"F0",X"F0",X"3C",X"F0",X"F0",
		X"F0",X"F0",X"0F",X"1E",X"3C",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"C3",X"87",X"0F",X"3C",X"F0",
		X"33",X"33",X"11",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"33",X"77",X"FF",
		X"00",X"FF",X"FF",X"FF",X"00",X"00",X"30",X"70",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"FF",X"EE",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"C0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"E0",X"F0",
		X"F0",X"10",X"00",X"30",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"EE",X"00",X"00",X"10",
		X"F0",X"10",X"F0",X"F0",X"F0",X"F0",X"70",X"80",X"F0",X"C0",X"10",X"E0",X"70",X"10",X"00",X"10",
		X"00",X"20",X"E0",X"D1",X"D1",X"D1",X"B3",X"80",X"00",X"00",X"00",X"10",X"70",X"30",X"30",X"00",
		X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",
		X"70",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"F0",X"EE",X"CC",X"CC",X"10",X"10",X"10",X"21",X"E1",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"78",X"1E",X"1E",
		X"F0",X"F0",X"E1",X"C3",X"E1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"F0",X"F0",X"3C",X"1E",X"0F",X"0F",X"F0",X"F0",X"78",X"1E",X"0F",X"0F",X"0F",X"C3",
		X"F0",X"70",X"F0",X"F0",X"F0",X"C3",X"0F",X"0F",X"70",X"00",X"F0",X"F0",X"F0",X"F0",X"78",X"0F",
		X"40",X"30",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"08",X"0F",X"0F",X"07",X"61",X"E1",X"C3",
		X"0F",X"07",X"00",X"80",X"C0",X"F0",X"F0",X"F0",X"0F",X"00",X"C0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"07",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"FF",X"0E",X"08",X"03",X"0F",X"07",X"00",X"EE",X"FF",
		X"0F",X"01",X"C0",X"3C",X"F0",X"E1",X"00",X"00",X"0C",X"78",X"3C",X"0F",X"F0",X"1C",X"00",X"CC",
		X"F0",X"3C",X"1E",X"0F",X"0F",X"0F",X"07",X"07",X"0F",X"0F",X"00",X"0E",X"0F",X"0F",X"00",X"88",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"C3",X"F0",X"0F",X"0F",X"0F",X"0F",X"C3",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"88",X"FF",X"FF",X"FF",X"FF",X"CC",X"FF",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0F",X"01",X"00",X"00",X"88",X"CC",X"0F",X"07",X"01",X"00",X"00",X"88",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"80",X"00",X"00",X"88",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"00",X"00",X"44",X"00",X"40",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"00",X"20",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"10",X"10",
		X"88",X"80",X"00",X"00",X"88",X"00",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"40",X"00",X"00",X"44",X"00",X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"20",X"00",X"00",X"22",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"10",X"00",X"00",X"11",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"C0",X"E8",X"E4",X"EC",X"E0",X"C0",X"00",X"00",X"10",X"30",X"30",X"30",X"10",X"00",X"00",
		X"00",X"E0",X"F4",X"F2",X"F6",X"F0",X"60",X"00",X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"70",X"F2",X"F1",X"F3",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",
		X"00",X"30",X"71",X"70",X"71",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C8",X"C8",X"C0",X"80",X"00",
		X"00",X"10",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E8",X"E4",X"EC",X"E0",X"C0",X"00",
		X"00",X"00",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"F4",X"F2",X"F6",X"F0",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"70",X"F2",X"F1",X"F3",X"70",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"80",X"C0",X"C8",X"C8",X"C0",X"80",X"00",X"00",X"30",X"71",X"70",X"71",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"E8",X"E4",X"EC",X"E0",X"C0",X"00",X"00",X"10",X"30",X"30",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"C0",X"E8",X"E4",X"EC",X"E0",X"00",X"00",X"00",X"10",X"30",X"30",X"30",X"10",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"E8",X"E4",X"EC",X"00",X"00",X"00",X"00",X"10",X"30",X"30",X"30",
		X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"E8",X"E4",X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"30",
		X"EC",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"30",
		X"E4",X"EC",X"E0",X"C0",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"E8",X"E4",X"EC",X"E0",X"C0",X"00",X"00",X"00",X"30",X"30",X"30",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C0",X"E8",X"E4",X"EC",X"E0",X"C0",X"00",X"00",X"10",X"30",X"30",X"30",X"10",X"00",X"00",X"00",
		X"80",X"F9",X"FE",X"F4",X"FE",X"FA",X"EC",X"C0",X"30",X"50",X"11",X"FD",X"91",X"30",X"C4",X"10",
		X"80",X"E8",X"F4",X"FF",X"F5",X"FE",X"FA",X"A0",X"00",X"64",X"91",X"98",X"33",X"D1",X"10",X"00",
		X"60",X"F6",X"F9",X"F6",X"FC",X"F5",X"FE",X"40",X"00",X"22",X"99",X"B3",X"B9",X"44",X"30",X"00",
		X"0C",X"02",X"01",X"11",X"F7",X"81",X"02",X"0C",X"03",X"04",X"18",X"58",X"78",X"38",X"04",X"03",
		X"0C",X"02",X"01",X"10",X"F8",X"89",X"02",X"0C",X"03",X"04",X"19",X"5D",X"7F",X"3B",X"04",X"03",
		X"0E",X"01",X"88",X"88",X"FC",X"CC",X"01",X"0E",X"01",X"02",X"04",X"26",X"37",X"15",X"02",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"80",X"08",X"00",X"00",
		X"0F",X"00",X"44",X"44",X"FE",X"EE",X"00",X"0F",X"00",X"01",X"02",X"13",X"13",X"02",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"40",X"C0",X"04",X"08",X"00",
		X"07",X"08",X"22",X"AA",X"FF",X"77",X"08",X"07",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"04",X"02",X"20",X"E0",X"02",X"04",X"08",
		X"03",X"04",X"19",X"5D",X"7F",X"3B",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"01",X"10",X"F8",X"89",X"02",X"0C",
		X"01",X"02",X"04",X"26",X"37",X"15",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"80",X"80",X"08",X"00",X"00",X"0E",X"01",X"88",X"88",X"FC",X"CC",X"01",X"0E",
		X"00",X"01",X"02",X"13",X"13",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"04",X"40",X"C0",X"04",X"08",X"00",X"0F",X"00",X"44",X"44",X"FE",X"EE",X"00",X"0F",
		X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"04",X"02",X"20",X"E0",X"02",X"04",X"08",X"07",X"08",X"22",X"AA",X"FF",X"77",X"08",X"07",
		X"00",X"00",X"88",X"F8",X"10",X"00",X"00",X"00",X"00",X"00",X"33",X"FF",X"DD",X"11",X"00",X"00",
		X"00",X"00",X"00",X"10",X"F8",X"88",X"00",X"00",X"00",X"00",X"11",X"DD",X"FF",X"33",X"00",X"00",
		X"00",X"0C",X"02",X"01",X"10",X"F8",X"89",X"02",X"00",X"03",X"04",X"19",X"5D",X"7F",X"3B",X"04",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"02",X"01",X"10",X"F8",X"89",X"00",X"00",X"03",X"04",X"19",X"5D",X"7F",X"3B",
		X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"02",X"01",X"10",X"F8",X"00",X"00",X"00",X"03",X"04",X"19",X"5D",X"7F",
		X"89",X"02",X"0C",X"00",X"00",X"00",X"00",X"00",X"3B",X"04",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"02",X"01",X"10",X"00",X"00",X"00",X"00",X"03",X"04",X"19",X"5D",
		X"F8",X"89",X"02",X"0C",X"00",X"00",X"00",X"00",X"7F",X"3B",X"04",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"03",X"04",X"19",
		X"10",X"F8",X"89",X"02",X"0C",X"00",X"00",X"00",X"5D",X"7F",X"3B",X"04",X"03",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"04",
		X"01",X"10",X"F8",X"89",X"02",X"0C",X"00",X"00",X"19",X"5D",X"7F",X"3B",X"04",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"02",X"01",X"10",X"F8",X"89",X"02",X"0C",X"00",X"04",X"19",X"5D",X"7F",X"3B",X"04",X"03",X"00",
		X"60",X"F7",X"EC",X"EA",X"F5",X"72",X"66",X"60",X"00",X"11",X"64",X"10",X"22",X"10",X"00",X"00",
		X"64",X"F9",X"F7",X"FE",X"FA",X"F7",X"FD",X"62",X"74",X"51",X"80",X"64",X"33",X"20",X"C4",X"00",
		X"62",X"F9",X"FA",X"F7",X"F4",X"FE",X"FB",X"64",X"88",X"20",X"A2",X"D8",X"00",X"F3",X"22",X"00",
		X"60",X"F6",X"F9",X"76",X"FC",X"F5",X"FE",X"62",X"33",X"40",X"BB",X"80",X"A8",X"44",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1E",X"1E",X"2C",X"2C",X"48",X"48",X"48",X"48",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"80",X"80",X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"3C",X"3C",
		X"C0",X"E0",X"68",X"68",X"68",X"48",X"48",X"48",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"3C",X"3C",X"68",X"68",X"68",X"48",X"C0",X"C0",X"F0",X"78",X"69",X"2D",X"2D",X"2D",X"0F",X"0F",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",
		X"F3",X"F3",X"F3",X"F3",X"71",X"70",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"48",X"48",X"68",X"2C",X"3C",X"3C",X"3C",X"3C",
		X"80",X"C0",X"C0",X"68",X"68",X"68",X"3C",X"3C",X"1E",X"0F",X"0F",X"2D",X"2D",X"69",X"78",X"F0",
		X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"3C",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",
		X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"30",X"70",X"71",X"F3",X"F3",X"F3",X"F3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"BB",X"30",X"30",X"33",X"33",X"30",X"30",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"30",X"30",X"33",X"33",X"B8",X"FC",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"FF",
		X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"00",
		X"AA",X"22",X"C5",X"E0",X"E0",X"C5",X"22",X"AA",X"88",X"55",X"75",X"F0",X"F0",X"75",X"55",X"88",
		X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"00",
		X"00",X"33",X"EE",X"CC",X"CC",X"EE",X"33",X"00",X"22",X"33",X"33",X"FF",X"FF",X"33",X"33",X"22",
		X"00",X"30",X"E0",X"C0",X"C0",X"E0",X"30",X"00",X"20",X"30",X"30",X"F0",X"F0",X"30",X"30",X"20",
		X"30",X"30",X"33",X"33",X"30",X"30",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"BB",X"30",X"30",X"33",X"33",X"30",X"30",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"30",X"30",X"33",X"33",X"B8",X"FC",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"FF",
		X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"0A",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"1C",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"09",X"00",X"80",X"08",X"09",X"0F",X"87",X"0C",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"1E",X"12",X"10",
		X"1E",X"1E",X"3C",X"78",X"F0",X"F0",X"F0",X"5A",X"09",X"00",X"80",X"08",X"09",X"0F",X"87",X"84",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"3C",X"78",X"3C",X"09",X"80",X"80",X"C0",X"C1",X"C3",X"C3",X"68",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"92",X"B0",X"80",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"2D",X"09",X"C0",X"C0",X"E0",X"F0",X"F0",X"B4",X"A4",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"C0",X"F0",X"F0",X"50",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"1E",X"09",X"C0",X"F0",X"F0",X"F0",X"F0",X"D2",X"58",
		X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0E",X"06",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"01",X"01",X"01",X"01",X"00",X"0B",X"0F",X"07",X"F6",X"ED",X"6B",X"6B",X"0F",X"0F",X"0F",X"0F",
		X"8E",X"0E",X"0E",X"0C",X"00",X"0E",X"1A",X"30",X"0B",X"0B",X"1C",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"0F",X"07",X"83",X"09",X"08",X"0C",X"87",X"0F",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"66",X"EE",X"88",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"1C",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"19",X"91",X"F3",X"7B",X"09",X"0F",X"87",X"0C",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"66",X"EE",X"88",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"1E",X"12",X"10",
		X"1E",X"1E",X"3C",X"78",X"F0",X"F0",X"F0",X"5A",X"19",X"91",X"F3",X"7B",X"09",X"0F",X"87",X"84",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"66",X"EE",X"88",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"3C",X"78",X"3C",X"19",X"91",X"F3",X"F3",X"C1",X"C3",X"C3",X"68",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"66",X"EE",X"88",X"0E",X"92",X"B0",X"80",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"2D",X"19",X"D1",X"F3",X"F1",X"F0",X"F0",X"B4",X"A4",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"00",X"00",X"02",X"03",X"01",X"0B",X"0F",X"07",X"0E",X"07",X"87",X"C3",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"66",X"EE",X"C0",X"F0",X"F0",X"50",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"1E",X"19",X"D1",X"F0",X"F0",X"F0",X"F0",X"D2",X"58",
		X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0E",X"06",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",
		X"01",X"01",X"01",X"01",X"00",X"0B",X"0F",X"07",X"F6",X"ED",X"6B",X"6B",X"0F",X"0F",X"0F",X"0F",
		X"8E",X"0E",X"0E",X"6E",X"EE",X"8E",X"1A",X"30",X"0B",X"0B",X"1C",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"0F",X"17",X"D3",X"59",X"7B",X"3F",X"87",X"0F",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"60",X"10",X"10",X"61",X"41",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"1E",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"09",X"00",X"80",X"08",X"09",X"0F",X"87",X"0C",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"60",X"10",X"10",X"61",X"41",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"1E",X"12",X"10",
		X"1E",X"1E",X"3C",X"78",X"F0",X"F0",X"F0",X"5A",X"09",X"00",X"80",X"08",X"09",X"0F",X"87",X"84",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"60",X"10",X"10",X"61",X"41",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"3C",X"78",X"3C",X"09",X"80",X"80",X"C0",X"C1",X"C3",X"C3",X"68",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"10",X"70",X"41",X"01",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"92",X"B0",X"80",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"2D",X"09",X"C0",X"C0",X"E0",X"F0",X"F0",X"B4",X"A4",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"10",X"70",X"41",X"01",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"C0",X"F0",X"F0",X"50",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"1E",X"09",X"C0",X"F0",X"F0",X"F0",X"F0",X"D2",X"58",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"60",X"10",X"10",X"61",X"41",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"C0",X"F0",X"F0",X"50",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"1E",X"09",X"C0",X"F0",X"F0",X"F0",X"F0",X"D2",X"58",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"60",X"10",X"10",X"61",X"41",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"92",X"B0",X"80",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"0F",X"0F",X"1E",X"3C",X"78",X"2D",X"09",X"C0",X"C0",X"E0",X"F0",X"F0",X"B4",X"A4",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"10",X"70",X"41",X"01",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"0F",X"03",X"01",
		X"1E",X"1E",X"1E",X"1E",X"1E",X"3C",X"78",X"3C",X"09",X"80",X"80",X"C0",X"C1",X"C3",X"C3",X"68",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"10",X"70",X"41",X"01",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"0D",X"0F",X"0F",X"1E",X"12",X"10",
		X"1E",X"1E",X"3C",X"78",X"F0",X"F0",X"F0",X"5A",X"09",X"00",X"80",X"08",X"09",X"0F",X"87",X"84",
		X"00",X"00",X"08",X"0C",X"04",X"8F",X"0F",X"0E",X"00",X"10",X"70",X"41",X"01",X"01",X"00",X"01",
		X"00",X"EE",X"FF",X"45",X"45",X"0B",X"0F",X"07",X"0E",X"07",X"8F",X"CB",X"4B",X"0F",X"0F",X"0F",
		X"0C",X"00",X"00",X"00",X"0E",X"1A",X"30",X"00",X"0B",X"0B",X"1E",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"09",X"00",X"80",X"08",X"09",X"0F",X"87",X"0C",
		X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0E",X"06",X"60",X"10",X"10",X"61",X"41",X"01",X"00",X"01",
		X"01",X"EF",X"EF",X"45",X"00",X"0B",X"0F",X"07",X"F6",X"ED",X"6B",X"6B",X"0F",X"0F",X"0F",X"0F",
		X"8E",X"0E",X"0E",X"0C",X"00",X"0E",X"1A",X"30",X"0B",X"0B",X"1C",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"0F",X"07",X"83",X"09",X"08",X"0C",X"87",X"0F",
		X"08",X"08",X"08",X"0C",X"0C",X"0C",X"0E",X"06",X"00",X"10",X"70",X"41",X"01",X"01",X"00",X"01",
		X"01",X"EF",X"EF",X"45",X"00",X"0B",X"0F",X"07",X"F6",X"ED",X"6B",X"6B",X"0F",X"0F",X"0F",X"0F",
		X"8E",X"0E",X"0E",X"0C",X"00",X"0E",X"1A",X"30",X"0B",X"0B",X"1C",X"3C",X"78",X"F0",X"E1",X"A1",
		X"1E",X"78",X"F0",X"E1",X"E1",X"F0",X"F0",X"B4",X"0F",X"07",X"83",X"09",X"08",X"0C",X"87",X"0F",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"30",X"F3",X"30",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"30",X"F3",X"30",X"00",X"00",X"0F",X"0F",X"08",
		X"73",X"73",X"73",X"00",X"05",X"2F",X"2F",X"22",X"F6",X"F6",X"F6",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",
		X"80",X"80",X"82",X"09",X"0F",X"87",X"86",X"C2",X"30",X"F3",X"30",X"00",X"00",X"0F",X"0F",X"08",
		X"75",X"75",X"75",X"00",X"05",X"2F",X"2F",X"22",X"FB",X"FB",X"FB",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"30",X"F3",X"30",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"FE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"B0",X"80",X"00",X"00",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"FE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"B0",X"80",X"00",X"00",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"30",X"F3",X"30",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"FE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"B0",X"80",X"00",X"00",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"FE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"B0",X"80",X"00",X"00",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"30",X"F3",X"30",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"FE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"B0",X"80",X"00",X"00",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",X"C8",
		X"88",X"88",X"8A",X"09",X"0F",X"87",X"86",X"C2",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"08",
		X"76",X"76",X"76",X"00",X"05",X"2F",X"2F",X"22",X"FD",X"FD",X"FD",X"C1",X"0C",X"1E",X"1C",X"50",
		X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"10",X"FE",X"88",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"F0",X"B0",X"80",X"00",X"00",X"62",X"40",X"C8",X"62",X"40",X"C8",X"62",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"11",X"00",X"80",X"50",X"00",X"22",X"00",X"00",X"00",X"00",X"20",X"44",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"54",X"80",X"00",X"11",X"00",X"00",X"00",X"00",X"40",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"20",X"00",X"89",X"73",X"1C",X"75",X"FB",X"00",X"00",X"00",X"95",X"C0",X"EC",X"C3",X"B2",
		X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"30",X"00",X"00",X"00",X"00",
		X"F9",X"EE",X"52",X"1A",X"00",X"00",X"00",X"00",X"E7",X"E8",X"06",X"48",X"15",X"80",X"00",X"00",
		X"00",X"44",X"00",X"00",X"10",X"00",X"00",X"40",X"00",X"22",X"00",X"01",X"00",X"41",X"01",X"03",
		X"00",X"00",X"0A",X"0B",X"0E",X"6C",X"F3",X"59",X"00",X"80",X"2C",X"0C",X"86",X"9F",X"C3",X"CF",
		X"00",X"00",X"00",X"22",X"80",X"00",X"44",X"00",X"03",X"10",X"01",X"00",X"80",X"00",X"00",X"00",
		X"F6",X"5E",X"2D",X"4B",X"02",X"88",X"00",X"00",X"46",X"86",X"8B",X"0E",X"08",X"04",X"00",X"80",
		X"00",X"00",X"28",X"08",X"04",X"48",X"2E",X"0C",X"00",X"10",X"01",X"00",X"24",X"03",X"03",X"07",
		X"11",X"03",X"0D",X"0F",X"4F",X"1E",X"C4",X"3E",X"0C",X"C5",X"0B",X"2B",X"9E",X"0F",X"43",X"8B",
		X"04",X"06",X"0E",X"84",X"00",X"88",X"80",X"00",X"07",X"01",X"02",X"07",X"23",X"16",X"01",X"00",
		X"2C",X"0E",X"B4",X"0F",X"07",X"2D",X"0E",X"CB",X"63",X"8B",X"4B",X"06",X"1F",X"9F",X"0D",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"55",X"77",X"00",X"77",X"44",X"77",X"00",X"44",X"44",X"CC",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"CC",X"44",X"CC",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"55",X"55",X"00",X"55",X"55",X"77",X"00",X"44",X"44",X"CC",X"00",X"CC",X"44",X"44",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"CC",X"44",X"CC",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"55",X"55",X"00",X"77",X"44",X"77",X"00",X"44",X"44",X"CC",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"CC",X"44",X"CC",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"44",X"77",X"44",X"00",X"77",X"44",X"77",X"00",X"88",X"CC",X"00",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"44",X"77",X"00",X"77",X"44",X"77",X"00",X"CC",X"44",X"CC",X"00",X"CC",X"44",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"44",X"77",X"44",X"00",X"77",X"44",X"00",X"00",X"88",X"CC",X"00",X"00",X"CC",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"77",X"44",X"77",X"00",X"00",X"00",X"CC",X"00",X"CC",X"44",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"22",X"3A",X"70",X"00",X"00",X"00",X"00",X"44",X"22",X"EA",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"3A",X"44",X"55",X"00",X"00",X"00",X"00",X"F0",X"EA",X"AA",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"44",X"3A",X"70",X"00",X"00",X"00",X"00",X"11",X"AA",X"EA",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"3A",X"22",X"11",X"00",X"00",X"00",X"00",X"F0",X"EA",X"22",X"44",X"00",X"00",X"00",X"00",
		X"F0",X"3B",X"63",X"E5",X"3B",X"30",X"88",X"41",X"38",X"33",X"3A",X"08",X"D1",X"3B",X"78",X"28",
		X"C4",X"40",X"40",X"E5",X"63",X"05",X"3B",X"C4",X"BE",X"E5",X"38",X"40",X"E4",X"C4",X"F0",X"41",
		X"30",X"5F",X"0A",X"3B",X"9C",X"E5",X"B2",X"89",X"3B",X"30",X"0C",X"B1",X"30",X"60",X"59",X"3B",
		X"20",X"FE",X"38",X"6B",X"5D",X"C4",X"40",X"88",X"6B",X"63",X"3B",X"3A",X"04",X"F6",X"19",X"78",
		X"0A",X"3B",X"00",X"21",X"1E",X"89",X"00",X"89",X"0C",X"B1",X"00",X"89",X"59",X"3B",X"00",X"89",
		X"38",X"00",X"89",X"89",X"40",X"00",X"89",X"89",X"3B",X"00",X"89",X"89",X"19",X"75",X"89",X"C8",
		X"E5",X"40",X"00",X"89",X"41",X"3B",X"60",X"61",X"08",X"38",X"14",X"29",X"28",X"F0",X"68",X"69",
		X"3A",X"F0",X"80",X"A8",X"08",X"00",X"C0",X"89",X"3A",X"00",X"88",X"E0",X"00",X"00",X"89",X"89",
		X"89",X"89",X"04",X"89",X"F0",X"F0",X"89",X"89",X"89",X"F0",X"89",X"89",X"F0",X"F0",X"89",X"4C",
		X"F0",X"A9",X"24",X"EA",X"A1",X"89",X"64",X"AB",X"E8",X"E1",X"2C",X"A3",X"89",X"89",X"6C",X"E3",
		X"F0",X"89",X"89",X"05",X"89",X"89",X"0C",X"45",X"89",X"89",X"F0",X"0D",X"89",X"89",X"44",X"4D",
		X"89",X"89",X"25",X"EB",X"89",X"F0",X"65",X"0E",X"89",X"89",X"2D",X"06",X"F0",X"E9",X"6D",X"46",
		X"4E",X"F0",X"AF",X"89",X"81",X"26",X"EF",X"50",X"F0",X"81",X"E7",X"18",X"07",X"2E",X"10",X"29",
		X"67",X"8F",X"89",X"89",X"86",X"CF",X"80",X"A8",X"6F",X"C7",X"89",X"C8",X"8E",X"A6",X"88",X"E0",
		X"0F",X"66",X"60",X"61",X"4F",X"27",X"21",X"89",X"47",X"6E",X"68",X"69",X"C1",X"2F",X"89",X"89",
		X"C6",X"AE",X"C0",X"89",X"CE",X"EE",X"89",X"89",X"C1",X"E6",X"89",X"89",X"87",X"A7",X"89",X"89",
		X"41",X"49",X"00",X"61",X"41",X"48",X"48",X"68",X"41",X"41",X"41",X"28",X"09",X"14",X"E0",X"BD",
		X"FF",X"27",X"08",X"01",X"68",X"21",X"00",X"49",X"49",X"63",X"A2",X"FF",X"28",X"41",X"40",X"09",
		X"08",X"FF",X"00",X"63",X"80",X"40",X"08",X"40",X"48",X"49",X"09",X"21",X"00",X"01",X"49",X"41",
		X"68",X"40",X"20",X"08",X"63",X"08",X"09",X"00",X"8A",X"69",X"41",X"A2",X"68",X"00",X"40",X"40",
		X"20",X"40",X"09",X"00",X"09",X"09",X"01",X"20",X"41",X"08",X"40",X"40",X"40",X"21",X"FF",X"41",
		X"20",X"49",X"49",X"09",X"09",X"08",X"08",X"01",X"41",X"40",X"09",X"40",X"40",X"A2",X"A2",X"FF",
		X"01",X"08",X"49",X"09",X"49",X"00",X"08",X"01",X"FF",X"4A",X"09",X"40",X"09",X"40",X"4A",X"FF",
		X"01",X"00",X"00",X"49",X"49",X"20",X"20",X"08",X"FF",X"40",X"40",X"09",X"09",X"41",X"41",X"07",
		X"00",X"49",X"FF",X"6B",X"20",X"41",X"09",X"40",X"40",X"09",X"49",X"00",X"41",X"08",X"40",X"20",
		X"41",X"2E",X"FF",X"40",X"40",X"40",X"09",X"41",X"09",X"00",X"49",X"20",X"01",X"20",X"49",X"09",
		X"09",X"2E",X"08",X"41",X"01",X"40",X"21",X"40",X"40",X"00",X"09",X"09",X"FF",X"20",X"08",X"01",
		X"FF",X"41",X"40",X"40",X"09",X"40",X"2E",X"FF",X"49",X"09",X"08",X"01",X"08",X"01",X"00",X"49",
		X"09",X"40",X"40",X"00",X"6B",X"FF",X"FF",X"20",X"08",X"01",X"01",X"40",X"00",X"49",X"49",X"41",
		X"40",X"09",X"49",X"09",X"41",X"C7",X"08",X"01",X"20",X"08",X"09",X"40",X"09",X"00",X"AF",X"FF",
		X"40",X"09",X"09",X"09",X"41",X"2E",X"08",X"01",X"20",X"08",X"41",X"40",X"09",X"00",X"AF",X"FF",
		X"40",X"40",X"00",X"49",X"FF",X"41",X"20",X"40",X"01",X"20",X"40",X"09",X"49",X"09",X"41",X"08",
		X"BA",X"DA",X"69",X"28",X"DA",X"DB",X"28",X"28",X"93",X"DA",X"69",X"69",X"DA",X"D3",X"28",X"28",
		X"F0",X"F0",X"28",X"F0",X"F0",X"F0",X"F0",X"F0",X"93",X"D2",X"69",X"DA",X"F0",X"F0",X"F0",X"F0",
		X"9A",X"D3",X"28",X"28",X"9A",X"F0",X"28",X"28",X"B2",X"9B",X"69",X"69",X"B2",X"F0",X"28",X"28",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"69",X"F0",X"F0",X"DA",X"9A",X"B2",X"D2",X"F0",X"69",X"F0",X"F0",
		X"F0",X"28",X"C3",X"0B",X"B3",X"28",X"23",X"0B",X"BA",X"69",X"0B",X"C3",X"FA",X"28",X"C4",X"23",
		X"28",X"69",X"23",X"02",X"28",X"8C",X"C3",X"0B",X"69",X"69",X"0B",X"23",X"28",X"02",X"0B",X"C3",
		X"FA",X"28",X"02",X"CC",X"28",X"28",X"02",X"02",X"F2",X"69",X"02",X"02",X"28",X"28",X"23",X"02",
		X"28",X"02",X"23",X"0B",X"69",X"23",X"02",X"8D",X"69",X"02",X"85",X"23",X"69",X"0B",X"02",X"02",
		X"02",X"02",X"0B",X"C3",X"23",X"02",X"AC",X"23",X"02",X"02",X"23",X"0B",X"0B",X"23",X"02",X"84",
		X"CD",X"23",X"0B",X"23",X"02",X"02",X"0B",X"C3",X"02",X"A4",X"C3",X"0B",X"02",X"02",X"23",X"0B",
		X"C3",X"0B",X"02",X"8C",X"23",X"0B",X"23",X"02",X"0B",X"C3",X"02",X"02",X"C5",X"23",X"0B",X"23",
		X"23",X"02",X"8C",X"23",X"C3",X"0B",X"02",X"8C",X"0B",X"23",X"8C",X"C4",X"0B",X"C3",X"02",X"02",
		X"02",X"02",X"23",X"0B",X"0B",X"23",X"8C",X"40",X"23",X"02",X"C5",X"23",X"C3",X"0B",X"02",X"40",
		X"8C",X"8D",X"40",X"40",X"02",X"02",X"40",X"40",X"02",X"8C",X"40",X"40",X"23",X"02",X"40",X"40",
		X"0B",X"C3",X"02",X"40",X"CC",X"23",X"0B",X"40",X"23",X"0B",X"23",X"40",X"8C",X"85",X"C3",X"40",
		X"0B",X"23",X"40",X"40",X"0B",X"C3",X"40",X"40",X"C3",X"0B",X"40",X"40",X"23",X"0B",X"40",X"A0",
		X"69",X"09",X"08",X"01",X"00",X"49",X"00",X"49",X"08",X"08",X"A2",X"FF",X"08",X"21",X"40",X"48",
		X"79",X"20",X"20",X"08",X"21",X"09",X"09",X"00",X"28",X"41",X"41",X"86",X"40",X"40",X"40",X"40",
		X"41",X"09",X"20",X"08",X"A0",X"20",X"09",X"00",X"48",X"40",X"41",X"86",X"00",X"08",X"40",X"40",
		X"08",X"01",X"01",X"20",X"00",X"49",X"49",X"09",X"A2",X"FF",X"FF",X"41",X"40",X"48",X"48",X"40",
		X"01",X"20",X"20",X"08",X"49",X"09",X"09",X"00",X"FF",X"41",X"41",X"99",X"48",X"40",X"40",X"40",
		X"08",X"01",X"01",X"20",X"00",X"49",X"49",X"09",X"19",X"FF",X"FF",X"41",X"40",X"48",X"48",X"40",
		X"08",X"01",X"01",X"20",X"00",X"49",X"49",X"09",X"19",X"FF",X"FF",X"41",X"40",X"48",X"48",X"40",
		X"20",X"08",X"08",X"01",X"09",X"00",X"00",X"49",X"41",X"99",X"C7",X"FF",X"40",X"40",X"40",X"48",
		X"08",X"01",X"01",X"20",X"00",X"49",X"49",X"09",X"C7",X"FF",X"FF",X"41",X"40",X"48",X"48",X"40",
		X"20",X"08",X"08",X"01",X"09",X"00",X"00",X"49",X"41",X"99",X"9C",X"FF",X"40",X"40",X"40",X"48",
		X"20",X"08",X"08",X"01",X"09",X"00",X"00",X"49",X"41",X"99",X"9C",X"FF",X"40",X"40",X"40",X"48",
		X"01",X"20",X"20",X"08",X"49",X"09",X"09",X"00",X"FF",X"41",X"41",X"5B",X"48",X"40",X"40",X"40",
		X"20",X"08",X"08",X"01",X"09",X"00",X"00",X"49",X"41",X"5B",X"19",X"FF",X"40",X"40",X"40",X"48",
		X"01",X"20",X"20",X"08",X"49",X"09",X"09",X"00",X"FF",X"41",X"41",X"5D",X"48",X"40",X"40",X"40",
		X"01",X"20",X"20",X"08",X"49",X"09",X"09",X"00",X"FF",X"41",X"41",X"5D",X"48",X"40",X"40",X"40",
		X"08",X"01",X"01",X"20",X"00",X"49",X"49",X"09",X"19",X"FF",X"FF",X"41",X"40",X"48",X"48",X"40");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
